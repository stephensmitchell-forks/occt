-- Created on: 1993-03-10
-- Created by: JCV
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RectangularTrimmedSurface from Geom inherits BoundedSurface from Geom

        ---Purpose : Describes a portion of a surface (a patch) limited
    	-- by two values of the u parameter in the u
    	-- parametric direction, and two values of the v
    	-- parameter in the v parametric direction. The
    	-- domain of the trimmed surface must be within the
    	-- domain of the surface being trimmed.
    	-- The trimmed surface is defined by:
    	-- - the basis surface, and
    	-- - the values (umin, umax) and (vmin, vmax)
    	--   which limit it in the u and v parametric directions.
    	--   The trimmed surface is built from a copy of the basis
    	-- surface. Therefore, when the basis surface is
    	-- modified the trimmed surface is not changed.
    	-- Consequently, the trimmed surface does not
    	-- necessarily have the same orientation as the basis surface.
	--  Warning:  The  case of surface   being trimmed is  periodic and
        --          parametrics values are outside the domain is possible.
    	--          But, domain of the  trimmed surface can be translated
    	--          by (n X) the period.

uses Ax1      from gp, 
     Ax2      from gp,
     Pnt      from gp,
     Trsf     from gp,
     GTrsf2d  from gp,
     Vec      from gp,
     Curve    from Geom, 
     Geometry from Geom,
     Shape    from GeomAbs,
     Surface  from Geom

raises ConstructionError   from Standard,
       RangeError          from Standard,
       NoSuchObject        from Standard,
       UndefinedDerivative from Geom,
       UndefinedValue      from Geom

is


  Create (S : Surface from Geom; 
          U1, U2, V1, V2 : Real; 
          USense, VSense : Boolean =  Standard_True)
     returns mutable RectangularTrimmedSurface
        ---Purpose :
        --  The U parametric direction of the surface is oriented from U1
        --  to U2. The V parametric direction of the surface is oriented 
        --  from V1 to V2.
        --  These two directions define the orientation of the surface 
        --  (normal). If the surface is not periodic USense and VSense are 
        --  not used for the construction. If the surface S is periodic in
        --  one direction USense and VSense give the available part of the
        --  surface. By default in this case the surface has the same
        --  orientation as the basis surface S.
        --  The returned surface is not closed and not periodic.
        --  ConstructionError   Raised if 
        --  S is not periodic in the UDirection and U1 or U2 are out of the 
        --  bounds of S.
        --  S is not periodic in the VDirection and V1 or V2 are out of the 
        --  bounds of S.
        --  U1 = U2 or V1 = V2

     raises ConstructionError;

  Create (S : Surface from Geom; 
          isUTrim, isVTrim : Boolean;
          U1, U2, V1, V2 : Real)
     returns mutable RectangularTrimmedSurface
        ---Purpose :
        --  The U parametric direction of the surface is oriented from U1
        --  to U2. The V parametric direction of the surface is oriented 
        --  from V1 to V2.
        --  These two directions define the orientation of the surface 
        --  (normal). By default in this case the surface has the same
        --  orientation as the basis surface S.
        --  isUTrim and isVTrim arguments determine, if it is necessary to
        --  trim S surface along corresponding direction.
        --  The returned surface is not closed and not periodic.
        --  ConstructionError   Raised if 
        --  S is not periodic in the UDirection and U1 or U2 are out of the 
        --  bounds of S.
        --  S is not periodic in the VDirection and V1 or V2 are out of the 
        --  bounds of S.
        --  U1 = U2 or V1 = V2

     raises ConstructionError;

     
  Create (S              : Surface from Geom; 
          Param1, Param2 : Real; 
          UTrim          : Boolean;
          Sense          : Boolean = Standard_True)
     returns mutable RectangularTrimmedSurface
        ---Purpose :
        --  The basis surface S is only trim in one parametric direction.
        --  If UTrim = True the surface is trimmed in the U parametric 
        --  direction else the surface is trimmed in the V parametric
        --  direction.
        --  In the considered parametric direction the resulting surface is
        --  oriented from Param1 to Param2. If S is periodic Sense gives the 
        --  available part of the surface. By default the trimmed surface has 
        --  the same orientation as the basis surface S in the considered 
        --  parametric direction (Sense = True).
        --  If the basis surface S is closed or periodic in the parametric
        --  direction opposite to the trimming direction the trimmed surface
        --  has the same characteristics as the surface S in this direction.
        -- Warnings :
        --  In this package the entities are not shared. 
        --  The RectangularTrimmedSurface is built with a copy of the 
        --  surface S. So when S is modified the RectangularTrimmedSurface
        --  is not modified
     raises ConstructionError;
        ---Purpose : Raised if 
        --  S is not periodic in the considered parametric direction and 
        --  Param1 or Param2 are out of the bounds of S.
        --  Param1 = Param2

    SetUTrim (me : mutable; U1, U2 : Real)
        ---Purpose : Sets boundaries of basisSurf in U1 and U2
        -- along U-direction.
        -- For periodic surface boundary values can be changed 
        -- algorithmically.
     raises ConstructionError;
        ---Purpose : Raised if 
        --  The BasisSurface is not periodic in the U-direction and U1 or U2
        --    are out of the bounds of the BasisSurface.
        --  U1 = U2

    SetVTrim (me : mutable; V1, V2 : Real)
        ---Purpose : Sets boundaries of basisSurf in V1 and V2
        -- along V-direction.
        -- For periodic surface boundary values can be changed 
        -- algorithmically.
     raises ConstructionError;
        ---Purpose : Raised if 
        --  The BasisSurface is not periodic in the V-direction and V1 or V2
        --    are out of the bounds of the BasisSurface.
        --  V1 = V2

    ForceTrim(me : mutable; 
              U1, U2, V1, V2 : Real; 
              UTrim, VTrim : Boolean = Standard_True);
      ---Purpose : For periodic surface this method changes
      -- (if it is necessary) U2 and V2, so that 0 < U2 - U1 < T and
      -- 0 < V2 - V1 < T (where T is the period).
      -- If surface is not periodic, boundaries do not chenge.
      -- After that it trims basisSurf in new boundaries.
        
  SetTrim (me : mutable; 
           U1, U2, V1, V2 : Real; 
           USense, VSense : Boolean = Standard_True)
        ---Purpose : Modifies this patch by changing the trim values
    	-- applied to the original surface
    	--        The u parametric direction of
    	--   this patch is oriented from U1 to U2. The v
    	--   parametric direction of this patch is oriented
    	--   from V1 to V2. USense and VSense are used
    	--   for the construction only if the surface is periodic
    	--   in the corresponding parametric direction, and
    	--   define the available part of the surface; by default
    	--   in this case, this patch has the same orientation
    	--   as the basis surface.
     raises ConstructionError;
        ---Purpose : Raised if 
        --  The BasisSurface is not periodic in the UDirection and U1 or U2
        --    are out of the bounds of the BasisSurface.
        --  The BasisSurface is not periodic in the VDirection and V1 or V2
        --    are out of the bounds of the BasisSurface.
        --  U1 = U2 or V1 = V2


  SetTrim (me : mutable; 
           Param1, Param2 : Real; 
           UTrim          : Boolean;
           Sense          : Boolean =  Standard_True)
        ---Purpose : Modifies this patch by changing the trim values
    	-- applied to the original surface
    	-- The basis surface is trimmed only in one parametric direction: if UTrim
    	--   is true, the surface is trimmed in the u parametric
    	--   direction; if it is false, it is trimmed in the v
    	--   parametric direction. In the "trimmed" direction,
    	--   this patch is oriented from Param1 to Param2. If
    	--   the basis surface is periodic in the "trimmed"
    	--   direction, Sense defines its available part. By
    	--   default in this case, this patch has the same
    	--   orientation as the basis surface in this parametric
    	--   direction. If the basis surface is closed or periodic
    	--   in the other parametric direction (i.e. not the
    	--   "trimmed" direction), this patch has the same
    	--  characteristics as the basis surface in that parametric direction. 
     raises ConstructionError;
        ---Purpose : Raised if 
        --  The BasisSurface is not periodic in the considered direction and
        --    Param1 or Param2 are out of the bounds of the BasisSurface.
        --  Param1 = Param2


  SetTrim (me : mutable; 
           U1, U2, V1, V2 : Real; 
	   UTrim, VTrim   : Boolean;
           USense, VSense : Boolean)
        ---Purpose :  General set trim,  to implement constructors and
        --         others set trim.
     raises ConstructionError
    is private;


  BasisSurface (me)   returns Surface from Geom;
        ---Purpose : Returns the Basis surface of <me>.


  UReverse (me : mutable);
    	---Purpose : Changes the orientation of this patch in the u 
    	-- parametric direction. The bounds of the surface are
    	-- not changed, but the given parametric direction is
    	-- reversed. Hence the orientation of the surface is reversed.
      

  UReversedParameter (me; U : Real) returns Real;
	---Purpose: Computes the u  parameter on the modified
    	-- surface, produced by when reversing its u 
    	-- parametric direction, for any point of u parameter U on this patch.
  
  VReverse (me : mutable);
    	---Purpose : Changes the orientation of this patch in the v
    	-- parametric direction. The bounds of the surface are
    	-- not changed, but the given parametric direction is
    	-- reversed. Hence the orientation of the surface is reversed.
       


  VReversedParameter (me; V : Real) returns Real;
    	---Purpose: Computes the v  parameter on the modified
    	-- surface, produced by when reversing its v 
    	-- parametric direction, for any point of v parameter V on this patch.
  
  Bounds (me; U1, U2, V1, V2 : out Real);
        ---Purpose : Returns the parametric bounds U1, U2, V1 and V2 of this patch.


  Continuity (me)  returns Shape from GeomAbs;
        ---Purpose : 
        --  Returns  the continuity of the surface : 
        --  C0 : only geometric continuity,
        --  C1 : continuity of the first derivative all along the Surface,
        --  C2 : continuity of the second derivative all along the Surface,
        --  C3 : continuity of the third derivative all along the Surface,
        --  CN : the order of continuity is infinite.


  IsUClosed (me)  returns Boolean;
    	---Purpose: Returns true if this patch is closed in the given parametric direction.

  IsVClosed (me)  returns Boolean;
    	---Purpose: Returns true if this patch is closed in the given parametric direction.

  IsCNu (me; N : Integer)  returns Boolean
        ---Purpose :
        --  Returns true if the order of derivation in the U parametric
        --  direction is N.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  IsCNv (me; N : Integer)  returns Boolean
        ---Purpose :
        --  Returns true if the order of derivation in the V parametric
        --  direction is N.
     raises RangeError;
        ---Purpose : Raised if N < 0.


  IsUPeriodic (me)  returns Boolean;
    	---Purpose: Returns true if this patch is periodic in the given
    	-- parametric direction.

  UPeriod (me)    returns Real from Standard
	---Purpose: Returns the period of this patch in the u 
    	-- parametric direction.
  raises
    	NoSuchObject from Standard
	---Purpose: raises if the surface is not uperiodic.
  is redefined;


  IsVPeriodic (me)  returns Boolean;
    	---Purpose:
    	-- Returns true if this patch is periodic in the given
    	-- parametric direction.
        
  VPeriod (me)    returns Real from Standard
	---Purpose: Returns the period of this patch in the v 
    	-- parametric direction.
  raises
    	NoSuchObject from Standard
	---Purpose: raises if the surface is not vperiodic.
  is redefined;



        ---Purpose : value and derivatives


  UIso (me; U : Real)  returns mutable Curve;
        ---Purpose : computes the U isoparametric curve.


  VIso (me; V : Real)   returns mutable Curve;
        ---Purpose : Computes the V isoparametric curve.


  D0 (me; U, V : Real; P : out Pnt)
     raises UndefinedValue;
        ---Purpose :
        --  Can be raised if the basis surface is an OffsetSurface.


  D1 (me; U, V : Real; P : out Pnt; D1U, D1V : out Vec)
        ---Purpose :
        --  The returned derivatives have the same orientation as the 
        --  derivatives of the basis surface even if the trimmed surface
        --  has not the same parametric orientation. 
    	--  Warning!  UndefinedDerivative  raised if the continuity of the surface is not C1.
     raises UndefinedDerivative;


  D2 (me; U, V : Real; P : out Pnt; D1U, D1V, D2U, D2V, D2UV : out Vec)
        --- Purpose :
        --  The returned derivatives have the same orientation as the 
        --  derivatives of the basis surface even if the trimmed surface
        --  has not the same parametric orientation.  
       -- Warning! UndefinedDerivative raised if the continuity of the surface is not C2.
     raises UndefinedDerivative;


  D3 (me; U, V : Real;  P : out Pnt; D1U, D1V, D2U, D2V, D2UV, 
      D3U, D3V, D3UUV, D3UVV : out Vec)
        --- Purposes : The returned derivatives have the same orientation as the 
        --  derivatives of the basis surface even if the trimmed surface
        --  has not the same parametric orientation. 
	        --  Warning UndefinedDerivative raised if the continuity of the surface is not C3.
     raises UndefinedDerivative;


  DN (me; U, V : Real; Nu, Nv : Integer)   returns Vec
        ---Purpose : The returned derivative has the same orientation as the 
        --  derivative of the basis surface even if the trimmed surface
        --  has not the same parametric orientation.
        --   Warning!  UndefinedDerivative raised if the continuity of the surface is not CNu in the U
        --  parametric direction and CNv in the V parametric direction.
        --  RangeError Raised if Nu + Nv < 1 or Nu < 0 or Nv < 0.    
     raises UndefinedDerivative,
  RangeError;



  Transform (me : mutable; T : Trsf);
    	---Purpose: Applies the transformation T to this patch.
    	-- Warning
    	-- As a consequence, the basis surface included in the
    	-- data structure of this patch is also modified.
    
  TransformParameters(me; U,V : in out Real; T : Trsf from gp)
	---Purpose: Computes the  parameters on the  transformed  surface for
	--          the transform of the point of parameters U,V on <me>.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are the new values of U,V after calling
	--          
	--          me->TranformParameters(U,V,T)
	--          
	--          This methods calls the basis surface method.
     is redefined;  

  ParametricTransformation(me; T : Trsf from gp) returns GTrsf2d from gp
	---Purpose: Returns a 2d transformation  used to find the  new
	--          parameters of a point on the transformed surface.
	--          
	--          me->Transformed(T)->Value(U',V')
	--          
	--          is the same point as
	--          
	--          me->Value(U,V).Transformed(T)
	--          
	--          Where U',V' are  obtained by transforming U,V with
	--          th 2d transformation returned by
	--          
	--          me->ParametricTransformation(T)
	--          
	--          This methods calls the basis surface method.
     is redefined;  

  Copy (me)  returns mutable like me;
    	---Purpose: Creates a new object which is a copy of this patch.
      
  GetTrimmedFlags(me; isUtrimmed,isVtrimmed : in out Boolean from Standard);
    	---Purpose: Allows to get <isutrimmed> and <isvtrimmed> members values.
      
fields

   basisSurf   : Surface from Geom;
   utrim1      : Real;
   vtrim1      : Real;
   utrim2      : Real;
   vtrim2      : Real;
   isutrimmed  : Boolean;
   isvtrimmed  : Boolean;

end;
