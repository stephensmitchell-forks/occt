-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AlgoTools2D from BOPTools 

      ---Purpose: 
      ---  The class contains handy static functions 
      ---  dealing with the topology  
      ---  This is the copy of the BOPTools_AlgoTools2D.cdl
uses 
    Vec  from gp, 
    Dir  from gp, 
    Vertex from TopoDS,
    Edge   from TopoDS, 
    Face   from TopoDS, 
     
    Curve from Geom2d,
    Curve from Geom, 
    ProjectedCurve from ProjLib

is   

    BuildPCurveForEdgeOnFace  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS); 
          ---Purpose: 
          --- Compute P-Curve for the edge <aE> on the face <aF> 
          ---
    EdgeTangent     (myclass;  
              anE  : Edge from TopoDS; 
              aT   : Real from Standard; 
              Tau  : out Vec  from gp) 
          returns  Boolean from Standard; 
          ---Purpose: 
          --- Compute tangent for the edge  <aE> [in 3D]  at parameter <aT> 
          ---
 
    PointOnSurface  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS;  
              aT:  Real from Standard; 
              U : out Real from Standard; 
              V : out Real from Standard); 
          ---Purpose: 
          --- Compute surface parameters <U,V> of the face <aF> 
          --- for  the point from the edge <aE> at parameter <aT>.   
          ---
    CurveOnSurface  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d; 
              aToler: out Real from Standard); 
          ---Purpose:  
          --- Get P-Curve <aC>  for the edge <aE> on surface <aF> . 
          --- If the P-Curve does not exist, build  it using Make2D(). 
          --- [aToler] - reached tolerance 
          ---
    CurveOnSurface  (myclass; 
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d; 
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard); 
                      
          ---Purpose: 
          --- Get P-Curve <aC>  for the edge <aE> on surface <aF> . 
          --- If the P-Curve does not exist, build  it using Make2D(). 
          --- [aFirst, aLast] - range of the P-Curve    
          --- [aToler] - reached tolerance 
          ---
    HasCurveOnSurface  (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d;
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard) 
          returns  Boolean from Standard; 
          ---Purpose:  
          --- Returns TRUE if the edge <aE>  has  P-Curve <aC>           
          --- on surface <aF> .   
          --- [aFirst, aLast] - range of the P-Curve    
          --- [aToler] - reached tolerance 
          --- If the P-Curve does not exist, aC.IsNull()=TRUE. 
          ---
    HasCurveOnSurface  (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS) 
          returns  Boolean from Standard;  
          ---Purpose:  
          --- Returns TRUE if the edge <aE>  has  P-Curve <aC>           
          --- on surface <aF> .   
          --- If the P-Curve does not exist, aC.IsNull()=TRUE. 
          ---
 
    AdjustPCurveOnFace  (myclass;    
              aF    :  Face from TopoDS; 
              C3D   :  Curve from Geom; 
              aC2D  :  Curve from Geom2d; 
              aC2DA : out Curve from Geom2d);                  
          ---Purpose:   
          --- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
          ---
    AdjustPCurveOnFace  (myclass;    
              aF    :  Face from TopoDS; 
              aT1   :  Real from Standard;   
              aT2   :  Real from Standard;   
              aC2D  :  Curve from Geom2d; 
              aC2DA : out Curve from Geom2d); 
          ---Purpose:   
          --- Adjust P-Curve <aC2D> (3D-curve <C3D>) on surface <aF> .  
          --- [aT1,  aT2] - range to adjust 
          ---
 
    IntermediatePoint (myclass; 
              aFirst: Real from Standard; 
              aLast : Real from Standard) 
          returns  Real from Standard; 
          ---Purpose:   
          --- Compute intermediate  value in  between [aFirst, aLast] . 
          ---
    IntermediatePoint        (myclass;  
              anE  : Edge from TopoDS) 
          returns  Real from Standard;
          ---Purpose:   
          --- Compute intermediate value of parameter for the edge <anE>. 
          ---
    BuildPCurveForEdgeOnPlane(myclass; 
              theE : Edge from TopoDS; 
              theF : Face from TopoDS);
 
    Make2D  (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d;
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard);            
          ---Purpose:   
          --- Make P-Curve <aC> for the edge <aE> on surface <aF> . 
          --- [aFirst, aLast] - range of the P-Curve    
          --- [aToler] - reached tolerance 
          --- 
          
    MakeCurveOnSurface        (myclass;  
              aE:  Edge from TopoDS; 
              aF:  Face from TopoDS; 
              aC    : out Curve from Geom2d;
              aFirst: out Real from Standard; 
              aLast : out Real from Standard; 
              aToler: out Real from Standard);             
          ---Purpose:   
          --- Same  as   Make2D() 
          ---
    MakePCurveOnFace  (myclass;    
              aF:  Face from TopoDS; 
              C3D   :     Curve from Geom; 
              aC    : out Curve from Geom2d; 
              aToler: out Real from Standard) ;   
          ---Purpose:   
          --- Make P-Curve <aC> for the 3D-curve <C3D> on surface <aF> . 
          --- [aToler] - reached tolerance 
          ---
    MakePCurveOnFace  (myclass;    
              aF:  Face from TopoDS; 
              C3D   :     Curve from Geom;  
              aT1   :  Real from Standard;   
              aT2   :  Real from Standard;      
              aC    : out Curve from Geom2d; 
              aToler: out Real from Standard) ;                  
          ---Purpose:   
          --- Make P-Curve <aC> for the 3D-curve <C3D> on surface <aF> .  
          --- [aT1,  aT2] - range to build    
          --- [aToler] - reached tolerance 
          ---
    MakePCurveOfType  (myclass;    
              PC  : ProjectedCurve from ProjLib; 
              aC  : out Curve from Geom2d);         
          ---Purpose:   
          --- Make empty  P-Curve <aC> of relevant to <PC> type  
          ---

 
 
 
 
 
 
 
--    RemovePCurveForEdgeOnFace  (myclass; 
--              aE:  Edge from TopoDS; 
--              aF:  Face from TopoDS); 
          ---Purpose: 
          --- Remove P-Curve of the edge <aE> on the face <aF> 
          ---
--    FaceNormal      (myclass; 
--              aF:  Face from TopoDS; 
--              U :  Real from Standard; 
--              V :  Real from Standard;  
--              aN: out Vec  from gp); 
          ---Purpose: 
          --- Compute normal for the face <aF> at parameters <U,V> 
          --- of the corresp. surface. 
          ---
--    TangentOnEdge    (myclass;  
--              aParm: Real from Standard; 
--              anE  : Edge from TopoDS;  
--              aTang: out Vec  from gp) 
--          returns  Boolean from Standard; 
--          ---Purpose:   
          --- Compute tangent for the edge <anE> at parameter <aParm>        
          ---
--    TangentOnEdge    (myclass;  
--              anE  : Edge from TopoDS;  
--              aDTang: out Dir  from gp) 
--          returns  Boolean from Standard;  
          ---Purpose:   
          --- Compute tangent for the edge <anE> at arbitrary intermediate parameter.        
          ---
--    TangentOnVertex  (myclass;  
--              aVF  : Vertex from TopoDS; 
--              aVL  : Vertex from TopoDS; 
--              anE  : Edge from TopoDS;  
--              aTang: out  Vec  from gp) 
--          returns  Boolean from Standard;  
          ---Purpose:   
          --- Compute tangent for the vertex point <aVF> for the edge <anE>. 
          --- <aVL> is opposite vertex of the edge        
          ---
--    EdgeBounds        (myclass; 
--              anE  : Edge from TopoDS;   
--              aFirst: out Real from Standard; 
--              aLast : out Real from Standard); 
          ---Purpose:   
          --- Returns parametric range for the edge <anE>. 
          ---

end AlgoTools2D;
