-- Created on: 2015-05-18
-- Created by: Sergey TELKOV
-- Copyright (c) 2015 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class IODevice from Storage inherits TShared from MMgt
    	---Purpose: Root any input output devices. A device define a way
    	-- to store or retrieve a data, for instance a file.

uses Position    from Storage,
     AsciiString from TCollection,
     OpenMode    from Storage,
     Error       from Storage,
     SeekMode    from Storage,
     ExtendedString from TCollection,
     SequenceOfAsciiString from TColStd,
     SequenceOfExtendedString from TColStd
     
raises StreamTypeMismatchError from Storage,
       StreamFormatError from Storage,
       StreamWriteError from Storage,
       StreamExtCharParityError from Storage
       
is
    Initialize;

    Delete( me : mutable ) is redefined;

    Name( me ) returns ExtendedString from TCollection is deferred;

    Open( me : mutable; aMode: OpenMode from Storage ) returns Error from Storage is deferred;

    OpenMode( me ) returns OpenMode from Storage;
    ---C++: inline

    IsEnd( me ) returns Boolean from Standard is deferred;
    ---Purpose: returns True if we are at end of the device data.

    Tell( me : mutable ) returns Position from Storage is deferred;
    ---Purpose: return position in the device. Return -1 upon error.

    Seek( me: mutable; aPos : Position from Storage; aMode: SeekMode from Storage = Storage_SMBegin )
    returns Boolean from Standard is deferred;
    ---Purpose: Set new absolute position within the stream
   
    Close(me : mutable) returns Boolean from Standard is deferred;

    CanRead(me) returns Boolean from Standard is deferred;

    CanWrite(me) returns Boolean from Standard is deferred;

    Read(me: mutable; aBuffer : Address from Standard;
                      aSize : Size from Standard)
    returns Size from Standard is deferred;

    Write(me: mutable; aBuffer : Address from Standard;
                       aSize : Size from Standard)
    returns Size from Standard is deferred;

    Signature(me) returns AsciiString from TCollection is deferred;

    Print(me; anOStream:  in out OStream from Standard)
    returns OStream from Standard is virtual;
    ---C++: return &
    ---C++: alias operator <<

    -- SERVICE

    ReadLine(me: mutable; aBuffer : in out CString from Standard; 
    	    	 aSize : Integer from Standard;
    	    	 anEndSymbol: Character from Standard);

    ReadLine(me: mutable; anEndSymbol: Character from Standard ) returns AsciiString from TCollection;


    WriteLine(me: mutable; aLine : CString from Standard);

    WriteLine(me: mutable; aLine : CString from Standard; anEndSymbol: Character from Standard);

    WriteLine(me: mutable; aLine : AsciiString from TCollection);

    WriteLine(me: mutable; aLine : AsciiString from TCollection; anEndSymbol: Character from Standard);

    -- PROTECTED

    SetOpenMode(me : mutable; aMode : OpenMode from Storage) is protected;
    ---C++: inline
    
fields

    myOpenMode : OpenMode from Storage;

end;
