-- Created on: 1992-02-03
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package Interface

    ---Purpose : defines a general frame for interface data
    --           used to manipulate results of normalized Interface outputs
    --           (i.e. files), also as a basis to define transfer operations
    --           (in other packages : see package Transfer)

uses LibCtl, TCollection, TColStd, MMgt, Standard, Dico, MoniTool, Message

is

    deferred class InterfaceModel;

    	-- --   Data Definitions   -- --

    class UndefinedContent;
    class ReportEntity;

    class EntityList;             -- for an (ordered) little list of Entities
    private class EntityCluster;  -- ancillary class for the former
    imported JaggedArray;    -- to turn arround limitation on Array(Array)

    	-- --   Auxiliary Classes (results, working data)   -- --

    class IntVal;
    class EntityIterator;

    class Graph;
    class GraphContent;
    class HGraph;
    class IntList;
    class BitMap;

    class Check;
    class CheckIterator;

    	-- --   General Services   -- --

    deferred class Protocol;         -- manages also Active Protocol
    deferred class GeneralModule;    -- (Shareds,Check,Copy,Trace)
    imported GeneralLib;

    class GTool;

    class ShareTool;
    class ShareFlags;
    class CheckTool;

    class CopyTool;
    deferred class CopyControl;
    class CopyMap;

    class Category;
    deferred class SignType;
    class SignLabel;

    class TypedValue;
    class Static;
    imported ValueSatisfies;
    -- (val : HAsciiString) returns Boolean,  see Satisfies from TypedValue
    imported ValueInterpret;
    -- (typval : TypedValue; hval : HAsciiString; native : Boolean)
    --   returns HAsciiString,  see Interpret from TypedValue
    imported StaticSatisfies;
    -- Function to be added to a Static for specific Satisfies

    imported Recognizer;  -- aimed to create Interface Entities

    	-- --   File Access (Read & Write)   -- --

    deferred class ReaderModule;
    imported ReaderLib;
    
    imported VectorOfFileParameter;
    class FileParameter;
    class ParamSet;          -- see also ParamList
    class ParamList;
    deferred class FileReaderData;
    deferred class FileReaderTool;

    class LineBuffer;
    class FloatWriter;

    class MSG;
    class STAT;

    	-- --   Enumerations   -- --

    enumeration ParamType is
    	ParamMisc, ParamInteger, ParamReal, ParamIdent, ParamVoid,   ParamText,
    	ParamEnum, ParamLogical, ParamSub,  ParamHexa,  ParamBinary;

    enumeration DataState is
    	StateOK, LoadWarning, LoadFail, DataWarning, DataFail,
    	StateUnloaded, StateUnknown;
    ---Purpose : validity state of anentity's content (see InterfaceModel)

    enumeration CheckStatus is
    	CheckOK, CheckWarning, CheckFail, CheckAny, CheckMessage, CheckNoFail;
    ---Purpose : Classifies checks
    --           OK : check is empty  Warning : Warning, no Fail   Fail : Fail
    --           Others to query :
    --           Any : any status   Message : Warning/Fail  NoFail : Warning/OK

    	-- --  Exceptions  -- --

    exception InterfaceError inherits Failure;
    exception InterfaceMismatch inherits InterfaceError;
    exception CheckFailure      inherits InterfaceError;

    	-- --  Instantiations  -- --

    private class  SequenceOfCheck  instantiates           -- for HSequence
    	 Sequence from TCollection (Check);
    private class HSequenceOfCheck  instantiates           -- Transient
    	HSequence from TCollection (Check,SequenceOfCheck);

    class Array1OfFileParameter instantiates               -- for ParamList :
        Array1 from TCollection    (FileParameter);
--    class HArray1OfFileParameter instantiates                           -- Array, Transient
--        HArray1 from TCollection   (FileParameter,Array1OfFileParameter);

    --  Useful Instantiations to define Data

    class  DataMapOfTransientInteger  instantiates  DataMap  from TCollection
    	(Transient, Integer,MapTransientHasher from TColStd);

    class  Array1OfHAsciiString instantiates   Array1  from TCollection
    	(HAsciiString from TCollection);

    class HArray1OfHAsciiString instantiates  HArray1  from TCollection
    	(HAsciiString from TCollection,Array1OfHAsciiString);

--  ==============IndexedMapOfAsciiString===================
class MapAsciiStringHasher;    -- instantiates MapHasher from TCollection;

class IndexedMapOfAsciiString instantiates IndexedMap  from TCollection(AsciiString from TCollection,MapAsciiStringHasher from Interface);

-- ==================================

end Interface;
