-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentStorageDriver from XmlLDrivers inherits StorageDriver from PCDM

uses
    AsciiString			from TCollection,
    ExtendedString		from TCollection,
    SequenceOfExtendedString	from TColStd,
    Document			from CDM,
    Document			from TDocStd,
    SequenceOfNamespaceDef	from XmlLDrivers,
    Element			from XmlObjMgt,
    SRelocationTable		from XmlObjMgt,
    ADriverTable		from XmlMDF,
    MessageDriver               from CDM,
    IODevice                    from Storage

is
    Create (theCopyright: ExtendedString from TCollection)
    	returns DocumentStorageDriver from XmlLDrivers;
    -- Constructor

    SchemaName(me) returns ExtendedString from TCollection is redefined virtual;
    -- pure virtual method definition

    Write	      (me: mutable;theDocument: Document       from CDM;
				   theDevice: IODevice from Storage)
	is redefined virtual;
    -- Write <aDocument> to the xml file <theFileName>

    WriteToDomDocument(me:mutable; theDocument: Document from CDM;
			           thePDoc    : out Element from XmlObjMgt;
   	    	    	    	   theDevice: IODevice from Storage)
	returns Boolean from Standard
	is virtual protected;

    MakeDocument      (me:mutable; theDocument: Document from CDM;
				   thePDoc    : out Element from XmlObjMgt)
	returns Integer from Standard
	is virtual protected;

    AddNamespace      (me:mutable; thePrefix, theURI: AsciiString)
	is protected;

    AttributeDrivers  (me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from XmlMDF
	is virtual; 
	
    WriteShapeSection (me:mutable; thePDoc    : out Element from XmlObjMgt) 
        returns Boolean from Standard
	is virtual protected; 
	
fields
    myDrivers   :	ADriverTable		 from XmlMDF is protected;
    mySeqOfNS	:	SequenceOfNamespaceDef	 from XmlLDrivers;
    myCopyright :       ExtendedString           from TCollection;
    myRelocTable:	SRelocationTable	 from XmlObjMgt  is protected;

end DocumentStorageDriver;
