-- Created on: 1998-03-27
-- Created by: Robert COUBLANC
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class Shape from StdSelect inherits PresentableObject from PrsMgr

	---Purpose: Presentable shape only for purpose of display for BRepOwner...

uses
    Projector             from Prs3d,
    Transformation        from Geom,
    Shape                 from TopoDS,
    PresentationManager3d from PrsMgr,
    Presentation          from Prs3d,
    Drawer                from Prs3d

is
    Create(Sh:Shape from TopoDS) returns mutable Shape from StdSelect;
    
    Compute(me:mutable;
    	        aPresentationManager: PresentationManager3d from PrsMgr;
                aPresentation: mutable Presentation from Prs3d;
                aMode: Integer from Standard = 0)
    is redefined static;
    
    Compute(me:mutable;
    	        aProjector: Projector from Prs3d;
                aPresentation: mutable Presentation from Prs3d)
    is redefined static private;     


    Compute(me            : mutable;
    	    aProjector    : Projector from Prs3d;
    	    aTrsf         : Transformation from Geom;
	    aPresentation : mutable Presentation from Prs3d)
    is redefined;
    	---Purpose: computes the presentation according to a point of view
    	--          given by <aProjector>. 
    	--          To be Used when the associated degenerated Presentations 
    	--          have been transformed by <aTrsf> which is not a Pure
    	--          Translation. The HLR Prs can't be deducted automatically
    	--          WARNING :<aTrsf> must be applied
    	--           to the object to display before computation  !!!

    Shape(me) returns Shape from TopoDS;
    	---C++: inline
    	---C++: return const&

    Shape(me:mutable;sh : Shape from TopoDS);
    	---C++: inline

    SetDrawer(me : mutable; aDrawer : Drawer from Prs3d);

fields
    mysh : Shape  from TopoDS;
    myDrawer : Drawer from Prs3d;
end Shape;
