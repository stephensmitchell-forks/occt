-- Created on: 1993-07-23
-- Created by: Martine LANGLOIS
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeBrepWithVoids from TopoDSToStep inherits
    Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Solid from TopoDS and BrepWithVoids from
    --          StepShape. All the topology and geometry comprised 
    --          into the shell or the solid are taken into account and
    --          translated.
  
uses Solid from TopoDS,
     BrepWithVoids from StepShape,
     FinderProcess_Handle from Transfer
          
raises NotDone from StdFail
     
is 

Create ( S  : Solid from TopoDS;
         FP : FinderProcess_Handle from Transfer)
        returns MakeBrepWithVoids;

Value (me) returns BrepWithVoids from StepShape
    raises NotDone
    is static;
    ---C++: return const&

fields

    theBrepWithVoids : BrepWithVoids from StepShape;

    	-- The solution from StepShape
    	
end MakeBrepWithVoids;


