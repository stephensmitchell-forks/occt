-- Created on: 1997-12-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private deferred class ReadWriter from PCDM inherits Transient from Standard

uses
    ExtendedString from TCollection,  
    AsciiString from TCollection, 
    Data from Storage, 
    Document from CDM, 
    MessageDriver from CDM,
    SequenceOfExtendedString from TColStd,  
    BaseDriver from Storage,  
    OpenMode from Storage, 
    SequenceOfReference from PCDM

is

    
    Version(me) returns AsciiString from TCollection
    is deferred;
    ---Purpose: returns PCDM_ReadWriter_1.
    
    WriteReferenceCounter(me; aData: Data from Storage; aDocument: Document from CDM)
    is deferred;
    
    WriteReferences(me; aData: Data from Storage; aDocument: Document from CDM; theReferencerFileName: ExtendedString from TCollection)
    is deferred;

    
    WriteExtensions(me; aData: Data from Storage; aDocument: Document from CDM)
    is deferred;

    
    WriteVersion(me; aData: Data from Storage; aDocument: Document from CDM)
    is deferred;

    
    ReadReferenceCounter(me; theFileName: ExtendedString from TCollection;   
			     theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard
    is deferred;

    ReadReferences(me; aFileName: ExtendedString from TCollection; theReferences: in out  SequenceOfReference from PCDM; theMsgDriver: MessageDriver from CDM)
    is deferred;

    ReadExtensions(me; aFileName: ExtendedString from TCollection; theExtensions: in out  SequenceOfExtendedString from TColStd; theMsgDriver: MessageDriver from CDM)
    is deferred;
    
    ReadDocumentVersion(me; aFileName: ExtendedString from TCollection; theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard
    is deferred;

---Category: commom methods


    Open(myclass; aDriver: in out BaseDriver from Storage; aFileName: ExtendedString from TCollection; anOpenMode: OpenMode from  Storage);
    
    Reader(myclass; aFileName: ExtendedString from TCollection)
    returns ReadWriter from PCDM;
    ---Purpose: returns the convenient Reader for a File.
    --          
    
    Writer(myclass)
    returns ReadWriter from PCDM;
    

    WriteFileFormat(myclass; aData: Data from Storage; aDocument: Document from CDM);
    
    FileFormat(myclass; aFileName: ExtendedString from TCollection)
    returns ExtendedString from TCollection;
    ---Purpose: tries  to get a format  in the  file.  returns an empty
    --          string if the file could not be read or does not have 
    --          a FileFormat information.

    FileFormat(myclass; theIStream: in out IStream from Standard; theData: out Data from Storage)
    returns ExtendedString from TCollection;

end ReadWriter from PCDM;
