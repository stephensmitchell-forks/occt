-- Created on: 1995-10-12
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepOffset 

	---Purpose: 

uses
    MMgt,
    Geom,
    TopoDS,
    TopAbs,	
    TCollection,
    TopTools,
    GeomAbs,
    BRepAlgo, 
    BOPAlgo, 
    BOPDS, 
    BOPTools

is
    enumeration Type is 
    	Concave, 
    	Convex, 
    	Tangent,
	FreeBoundary,
	Other
    end Type;
    
    enumeration Mode is 
    	Skin,
    	Pipe,
    	RectoVerso 
    end Mode;
---Purpose:
-- Lists the offset modes. These are the following:
-- - BRepOffset_Skin which describes the offset along
--   the surface of a solid, used to obtain a manifold topological space,
-- - BRepOffset_Pipe which describes the offset of a
--   curve, used to obtain a pre-surface,
-- - BRepOffset_RectoVerso which describes the offset
--   of a given surface shell along both sides of the surface.
        
    enumeration Status is 
	---Purpose: status of an offset face
	--          Good : 
	--          Reversed : e.g. Offset > Radius of a cylinder
	--          Degenerated : e.g. Offset = Radius of a cylinder
	--          Unknown : e.g. for a Beziersurf
    	Good,
	Reversed,
	Degenerated,
    	Unknown
    end Status;
    	    
    enumeration Error is
        NoError,		    	
	OffsetSurfaceFailed,
	UnCorrectClosingFace,
        ExtentFaceFailed,
	RadiusEqualOffset,
	UnknownError
    end Error;
    
    class MakeOffset;
    class MakeOffsetOld;
    	
    --class Loop;
    
    class Inter3d;
    
    class Inter2d;
    
    class Offset;

    class Analyse;

    class MakeLoops;
    
    class Tool;

    --class Image;
    
    --class AsDes;


    class Interval;
   
    class ListOfInterval instantiates 
    	List from TCollection  (Interval from BRepOffset);
    
    class DataMapOfShapeListOfInterval  instantiates
    	DataMap from TCollection(Shape           from TopoDS,
	    	    	    	 ListOfInterval  from BRepOffset,
				 ShapeMapHasher  from TopTools );   
    
    class DataMapOfShapeOffset instantiates
    	DataMap from TCollection(Shape           from TopoDS,
	    	    	    	 Offset          from BRepOffset,
				 ShapeMapHasher  from TopTools );   
				 
    class DataMapOfShapeMapOfShape instantiates
	DataMap from TCollection(Shape           from TopoDS,
	    	    	    	 MapOfShape      from TopTools,
				 ShapeMapHasher  from TopTools);     

  
    Surface( Surface : in  Surface from Geom;
    	     Offset  : in  Real    from Standard;
    	     Status  : out Status  from BRepOffset)
	---Purpose: returns   the  Offset  surface  computed from  the
	--          surface <Surface> at an OffsetDistance <Offset>.
	--          
	--          If possible, this method returns  the real type of
	--          the surface ( e.g. An Offset of a plane is a plane).
	--          
	--          If  no particular  case  is detected, the returned
	--          surface will have the Type Geom_OffsetSurface.
    returns Surface from Geom;

end BRepOffset;
