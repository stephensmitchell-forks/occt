-- Created on: 1992-02-04
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TransferInput  from Transfer

    ---Purpose : A TransferInput is a Tool which fills an InterfaceModel with
    --           the result of the Transfer of CasCade Objects, once determined
    --           The Result comes from a TransferProcess, either from
    --           Transient (the Complete Result is considered, it must contain
    --           only Transient Objects)

uses InterfaceModel, EntityIterator, Protocol from Interface,
     TransferIterator, TransientProcess_Handle, FinderProcess_Handle

raises TransferFailure

is

    Create returns TransferInput;
    ---Purpose : Creates a TransferInput ready to use

    Entities (me; list : in out TransferIterator) returns EntityIterator
    ---Purpose : Takes the transient items stored in a TransferIterator
    	raises TransferFailure;
    --           Error if one of the Resulting Objects is defined not Transient


    FillModel (me; proc   : TransientProcess_Handle;
    	    	   amodel : mutable InterfaceModel)
    ---Purpose : Fills an InterfaceModel with the Complete Result of a Transfer
    --           stored in a TransientProcess (Starting Objects are Transient)
    --           The complete result is exactly added to the model
    	raises TransferFailure;
    --           Error if one of the Resulting Objects is defined not Transient

    FillModel (me; proc   : TransientProcess_Handle;
    	    	   amodel : mutable InterfaceModel;
		   proto  : Protocol from Interface;
		   roots  : Boolean = Standard_True)
    ---Purpose : Fills an InterfaceModel with results of the Transfer recorded
    --           in a TransientProcess (Starting Objects are Transient) :
    --           Root Result if <roots> is True (Default), Complete Result else
    --           The entities added to the model are determined from the result
    --           by by adding the referenced entities
    	raises TransferFailure;
    --           Error if one of the Resulting Objects is defined not Transient


    FillModel (me; proc   : FinderProcess_Handle;
    	    	   amodel : mutable InterfaceModel)
    ---Purpose : Fills an InterfaceModel with the Complete Result of a Transfer
    --           stored in a TransientProcess (Starting Objects are Transient)
    --           The complete result is exactly added to the model
    	raises TransferFailure;
    --           Error if one of the Resulting Objects is defined not Transient

    FillModel (me; proc   : FinderProcess_Handle;
    	    	   amodel : mutable InterfaceModel;
		   proto  : Protocol from Interface;
		   roots  : Boolean = Standard_True)
    ---Purpose : Fills an InterfaceModel with results of the Transfer recorded
    --           in a TransientProcess (Starting Objects are Transient) :
    --           Root Result if <roots> is True (Default), Complete Result else
    --           The entities added to the model are determined from the result
    --           by by adding the referenced entities
    	raises TransferFailure;
    --           Error if one of the Resulting Objects is defined not Transient

end TransferInput;
