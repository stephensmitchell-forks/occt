-- Created on: 1994-06-16
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package HeaderSection 

uses


	TCollection, TColStd, StepData, Interface, MMgt

is



class Protocol;


class FileName;
class FileDescription;
class FileSchema;

imported HeaderRecognizer;

--class Array1OfHAsciiString instantiates Array1(HAsciiString);
--class HArray1OfHAsciiString instantiates HArray1(HAsciiString,Array1OfHAsciiString from HeaderSection);
-- already instantiated in package Interface

	Protocol returns Protocol from HeaderSection;
	---Purpose : creates a Protocol

end HeaderSection;

