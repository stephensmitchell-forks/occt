-- Created on: 1998-06-03
-- Created by: data exchange team
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package ShapeFix 

  ---Purpose:  This package provides algorithms for fixing
  -- problematic (violating Open CASCADE requirements) shapes.
  -- Tools from package ShapeAnalysis are used for detecting the problems. The
  -- detecting and fixing is done taking in account various
  -- criteria implemented in BRepCheck package. 
  -- Each class of package ShapeFix deals with one
	-- certain type of shapes or with some family of problems.

uses

    gp,
    Geom,
    Geom2d,
    Geom2dAPI,
    GeomAbs,
    Adaptor3d,
    TCollection,
    TColStd,
    TopAbs,
    TopLoc,
    TopoDS, 
    TopTools,
    Message,
    ShapeExtend,
    ShapeAnalysis,
    ShapeConstruct,
    ShapeBuild,
    Bnd

is

    -- classes
    class Root;    

    class EdgeProjAux;

    class Edge;
    	---Purpose: Fixing different problems on edge
	
    class Wire;
      ---Purpose: Fixing different problems with wires

    class Face;
    	---Purpose: Fixing problems with face (orientation of wires and wrong wires)
	  
    class FixSmallFace;
      ---Purpose: Fixing face with small size

    class WireVertex;
    	---Purpose: Fixing disconnected edges in the wire

    class Wireframe;
      ---Purpose: Provides methods to fix wireframe of shape
    
    class FreeBounds;
      ---Purpose: Fixing free bounds of the shape (connecting open wires)

    class FaceConnect;
      ---Purpose: Rebuilds connectivity between faces in shell
	
    class Shell;
    	---Purpose: Fixing orientation of faces in shell

    class Solid;
      ---Purpose: Creating solid from shell and orienting it to have finite volume
	
    class ShapeTolerance;
    	---Purpose: Modifying shape tolerances

    class Shape;
    	---Purpose: Fixing problem of shape. 

    class EdgeConnect;
        ---Purpose: Rebuilds edges to connect with new vertices, was moved from ShapeBuild

    class ComposeShell;
    	---Purpose: Splits a (pseudo)face onto grid of faces (shell)

    class SplitCommonVertex;
    	---Purpose: Splits vertex which is common for two wires
      --          (for writing into STEP)

    class WireSegment;
    	---Purpose: Auxiliary class (data storage) for ComposeShell
	
    class IntersectionTool;
    	---Purpose: Tool for fixing selfintersecting wire
      --          and intersecting wires
	
    class SplitTool;
    	---Purpose: Tool for splitting and cutting edges; incudes methods
      --          used in OverlappingTool and IntersectionTool
	
    class SequenceOfWireSegment instantiates Sequence from TCollection
    	(WireSegment from ShapeFix);
    
    class DataMapOfShapeBox2d instantiates DataMap from TCollection                           
    	(Shape from TopoDS, Box2d from Bnd, ShapeMapHasher from TopTools);


    SameParameter (shape       : Shape from TopoDS;
                   enforce     : Boolean;
                   preci       : Real = 0.0;
                   theProgress : ProgressIndicator from Message = 0)
    returns Boolean;
    	---Purpose : Runs SameParameter from BRepLib with these adaptations :
    	--           <enforce> forces computations, else they are made only on
    	--             Edges with flag SameParameter false
    	--           <preci>, if not precised, is taken for each EDge as its own
    	--           Tolerance
    	--           Returns True when done, False if an exception has been raised
    	--           In case of exception anyway, as many edges as possible have
    	--           been processed. The passed progress indicator allows user
    	--           to consult the current progress stage and abort algorithm
    	--           if needed.

    EncodeRegularity (shape: Shape from TopoDS; tolang: Real = 1.0e-10);
    	---Purpose : Runs EncodeRegularity from BRepLib taking into account
      --           shared components of assemblies, so that each component
      --           is processed only once

    RemoveSmallEdges (shape: in out Shape from TopoDS; Tolerance: Real; context: in out ReShape from ShapeBuild) 
    	returns Shape from TopoDS;
      ---Purpose: Removes edges which are less than given tolerance from shape
      --          with help of ShapeFix_Wire::FixSmall()

    FixVertexPosition(theshape: in out Shape from TopoDS;
		      theTolerance: Real; 
    	    	      thecontext: ReShape from ShapeBuild) returns Boolean;
      ---Purpose: Fix position of the vertices having tolerance more tnan specified one.;       
    	 
    LeastEdgeSize(theshape: in out Shape from TopoDS) returns Real;
      ---Purpose: Calculate size of least edge;       

    RefineFace (theF        :        Face  from TopoDS;
                theNewShape : in out Shape from TopoDS;
                flForce : Boolean from Standard = Standard_False;
                flDoNotSplit : Boolean from Standard = Standard_True);
    ---Purpose: It is created for fixing faces with 
    --          BRepCheck_OutOfSurfaceBoundary status.
    --          If source face is based on not RectangularTrimmed
    --          surface and after this method calling it should be 
    --          based on RectangularTrimmed surface (for successfull
    --          fixing), then fixing will be executed if and only if
    --          flForce == Standard_True.
    --          If it is necessary to do splitting, flForce allows to
    --          ignore periodic of source surface, which theF based on.
    --          flDoNotSplit forbids to split principial.
		
    ReTrimmedFace(theF        : in out Face       from TopoDS;
                  theNewRTSurf: RectangularTrimmedSurface from Geom)
                  
    ---Purpose:    Replace the surface in theF with theNewRTSurf.
    is private;
    
    SplittingFace(theF        :        Face  from TopoDS;
                  theNewShape : in out Shape from TopoDS;
                  theS  : Surface from Geom;
                  theDeltaBU2, theDeltaBV2,
                  theUFf, theVFf,
                  theUReminder, theVReminder : Real from Standard;
                  isSplitByU, isSplitByV : Boolean from Standard)
                  
    ---Purpose:    Make split.
    is private;
      
end ShapeFix;
