-- Created on: 2004-01-09
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DimTolTool from XCAFDoc inherits Attribute from TDF

	---Purpose: Provides tools to store and retrieve attributes (colors)
	--          of TopoDS_Shape in and from TDocStd_Document
	--          A Document is intended to hold different 
	--          attributes of ONE shape and it's sub-shapes.
	--          Attribute containing DimTol section of DECAF document.
	--          Provide tools for management of DimTol section of document.
uses
    Shape from TopoDS,
    Label from TDF,
    LabelSequence from TDF,
    Document from TDocStd,
    ShapeTool from XCAFDoc,
    GeomTolerance from XCAFDoc,
    Datum from XCAFDoc,
    Dimension from XCAFDoc,
    RelocationTable from TDF,
    HArray1OfReal from TColStd,
    HAsciiString from TCollection

is
    Create returns DimTolTool from XCAFDoc;

    Set (myclass; L : Label from TDF) returns DimTolTool from XCAFDoc;
    	---Purpose: Creates (if not exist) DimTolTool.
    
    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;

    
    
    ---API: General structure
    
    BaseLabel(me) returns Label from TDF;
    	---Purpose: returns the label under which colors are stored
    
    ShapeTool (me: mutable) returns ShapeTool from XCAFDoc;
    	---Purpose: Returns internal XCAFDoc_ShapeTool tool
	---C++: return const &



    -- Methods for Dimension:

    IsDimension (me; theLab: Label from TDF) returns Boolean;
    	---Purpose: Returns True if label belongs to a dimtoltable and
        --          is a Dimension definition 

    GetDimensionLabels (me; theLabels: out LabelSequence from TDF);
    	---Purpose: Returns a sequence of Dimensions labels currently stored 
        --          in the DGTtable


    SetDimension (me; theFirstL: Label from TDF;
                   theSecondL: Label from TDF;
		   theDimTolL: Label from TDF);
    	---Purpose: Sets a link with GUID

    SetDimension (me; theL: Label from TDF;
		   theDimTolL: Label from TDF);
    	---Purpose: Sets a link with GUID

    GetRefDimensionLabels (me; theShapeL: Label from TDF; theDimensions: out LabelSequence from TDF) 
    returns Boolean;
    	---Purpose: Returns all Dimension labels defined for label ShapeL

    AddDimension (me : mutable)
    returns Label from TDF;
    	---Purpose: Adds a dimension definition to a DGTtable and returns its label



    -- Methods for GeomTolerance:

    IsGeomTolerance (me; theLab: Label from TDF) returns Boolean;
    	---Purpose: Returns True if label belongs to a dimtoltable and
        --          is a DimTol definition 

    GetGeomToleranceLabels (me; theLabels: out LabelSequence from TDF);
    	---Purpose: Returns a sequence of Tolerance labels currently stored 
        --          in the DGTtable

    SetGeomTolerance (me; theL: Label from TDF;
		   theDimTolL: Label from TDF);
    	---Purpose: Sets a link with GUID

    GetRefGeomToleranceLabels (me; theShapeL: Label from TDF; theDimTols: out LabelSequence from TDF) 
    returns Boolean;
    	---Purpose: Returns all GeomTolerance labels defined for label ShapeL

    AddGeomTolerance (me : mutable)
    returns Label from TDF;
    	---Purpose: Adds a GeomTolerance definition to a DGTtable and returns its label



    -- Methods for DimTol:

    IsDimTol (me; lab: Label from TDF) returns Boolean;
    	---Purpose: Returns True if label belongs to a dimtoltable and
        --          is a DimTol definition 
    
    GetDimTolLabels (me; Labels: out LabelSequence from TDF);
    	---Purpose: Returns a sequence of D&GTs currently stored 
        --          in the DGTtable
    
    FindDimTol (me; kind : Integer from Standard; aVal : HArray1OfReal from TColStd;
    	    	    aName : HAsciiString from TCollection;
		    aDescription : HAsciiString from TCollection;
                    lab: out Label from TDF)
    returns Boolean;
    	---Purpose: Finds a dimtol definition in a DGTtable and returns
	--          its label if found
    	--          Returns False if dimtol is not found in DGTtable 
    
    FindDimTol (me; kind : Integer from Standard; aVal : HArray1OfReal from TColStd;
    	    	    aName : HAsciiString from TCollection;
    	    	    aDescription : HAsciiString from TCollection)
    returns Label from TDF;
    	---Purpose: Finds a dimtol definition in a DGTtable and returns
	--          its label if found (or Null label else)
    
    AddDimTol (me; kind : Integer from Standard;
    	    	   aVal : HArray1OfReal from TColStd;
    	    	   aName : HAsciiString from TCollection;
    	    	   aDescription : HAsciiString from TCollection)
    returns Label from TDF;
    	---Purpose: Adds a dimtol definition to a DGTtable and returns its label

    SetDimTol (me; L: Label from TDF;
		   DimTolL: Label from TDF);
    	---Purpose: Sets a link with GUID
    
    SetDimTol (me; L: Label from TDF; kind : Integer from Standard;
    	    	   aVal : HArray1OfReal from TColStd;
    	    	   aName : HAsciiString from TCollection;
    	    	   aDescription : HAsciiString from TCollection)
    returns Label from TDF;
    	---Purpose: Sets a link with GUID
    	--          Adds a DimTol as necessary
    
    GetRefShapeLabel (me; theDimTolL: Label from TDF; theShapeL: out LabelSequence from TDF) 
    returns Boolean;
    	---Purpose: Returns ShapeL defined for label DimTolL
	--          Returns False if the DimTolL is not in DGTtable

    GetRefDGTLabels (me; theShapeL: Label from TDF; theDimTols: out LabelSequence from TDF) 
    returns Boolean;
    	---Purpose: Returns all DimTol labels defined for label ShapeL

    GetDimTol (me; DimTolL: Label from TDF; kind : out Integer from Standard;
    	    	   aVal : out HArray1OfReal from TColStd;
    	    	   aName : out HAsciiString from TCollection;
    	    	   aDescription : out HAsciiString from TCollection) returns Boolean;
        ---Purpose: Returns dimtol assigned to <DimTolL>
    	--          Returns False if no such dimtol is assigned
    

    -- Methods for Datum:

    IsDatum (me; theLab: Label from TDF) returns Boolean;
    	---Purpose: Returns True if label belongs to a dimtoltable and
        --          is a Datum definition 
    
    GetDatumLabels (me; theLabels: out LabelSequence from TDF);
    	---Purpose: Returns a sequence of Datum labels currently stored 
        --          in the DGTtable
   
    FindDatum (me; aName : HAsciiString from TCollection;
		   aDescription : HAsciiString from TCollection;
		   anIdentification : HAsciiString from TCollection;
                   lab: out Label from TDF)
    returns Boolean;
    	---Purpose: Finds a datum and returns its label if found
    
    AddDatum (me; aName : HAsciiString from TCollection;
    	    	  aDescription : HAsciiString from TCollection;
    	    	  anIdentification : HAsciiString from TCollection)
    returns Label from TDF;
    	---Purpose: Adds a datum definition to a DGTtable and returns its label

    AddDatum (me : mutable)
    returns Label from TDF;
    	---Purpose: Adds a datum definition to a DGTtable and returns its label

    SetDatum (me; theL: Label from TDF;
		  theDatumL: Label from TDF);
    	---Purpose: Sets a link with GUID
    
    SetDatum (me; L: Label from TDF; TolerL: Label from TDF;
    	    	  aName : HAsciiString from TCollection;
    	    	  aDescription : HAsciiString from TCollection;
    	    	  anIdentification : HAsciiString from TCollection);
    	---Purpose: Sets a link with GUID for Datum
    	--          Adds a Datum as necessary
	--          Sets connection between Datum and Tolerance

    SetDatumToGeomTol (me; theL: Label from TDF; theTolerL: Label from TDF);
    	---Purpose: Sets a link with GUID for Datum
	--          Sets connection between Datum and Tolerance

    
    GetDatum (me; DatumL: Label from TDF;
    	    	  aName : out HAsciiString from TCollection;
    	    	  aDescription : out HAsciiString from TCollection;
                  anIdentification : out HAsciiString from TCollection) returns Boolean;
        ---Purpose: Returns datum assigned to <DatumL>
    	--          Returns False if no such datum is assigned
    
    GetDatumOfTolerLabels (me; theDimTolL: Label from TDF; theDatums: out LabelSequence from TDF) 
    returns Boolean;
    	---Purpose: Returns all Datum labels defined for label DimTolL

    GetTolerOfDatumLabels (me; theDatumL: Label from TDF; theTols: out LabelSequence from TDF) 
    returns Boolean;
    	---Purpose: Returns all GeomToleranses labels defined for label DatumL

    GetRefDatumLabel (me; theShapeL: Label from TDF; theDatum: out Label from TDF) 
    returns Boolean;
    	---Purpose: Returns Datum label defined for label ShapeL

    GetRefDatum (me; theShape: Shape from TopoDS; theDatum: out Datum from XCAFDoc) 
    returns Boolean;
    	---Purpose: Returns Datum label defined for label Shape

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

fields

    myShapeTool: ShapeTool from XCAFDoc;
    
end DimTolTool;
