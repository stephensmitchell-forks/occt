-- Created on: 1992-09-30
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class QuadricTool from IntSurf

	---Purpose: This class provides a tool on a quadric that can be
	--          used to instantiates the Walking algorithmes (see
	--          package IntWalk) with a Quadric from IntSurf
	--          as implicit surface.

uses Quadric from IntSurf,
     Vec     from gp,
     Pnt     from gp

is

    Value(myclass; Quad: Quadric from IntSurf;
          X, Y, Z: Real from Standard)
	  
    	---Purpose: Returns the value of the function.
    
    	returns Real from Standard;
	
	---C++: inline
    
    
    Gradient(myclass; Quad: Quadric from IntSurf;
             X, Y, Z: Real from Standard ; V : out Vec from gp);
	     
    	---Purpose: Returns the gradient of the function.

	---C++: inline
    


    ValueAndGradient(myclass; Quad: Quadric from IntSurf;
                     X, Y, Z: Real from Standard;
                     Val: out Real from Standard;
    	    	     Grad: out Vec from gp;
		     D1U_ISurf, D1V_ISurf: out Vec from gp);
		     
    	---Purpose: Returns the value and the gradient.

    D2(myclass; Quad:  Quadric from IntSurf;
                Point: Pnt from gp;
    	    	D1U:   out Vec from gp;
    	    	D1V:   out Vec from gp;
    	    	D2U:   out Vec from gp;
    	    	D2V:   out Vec from gp;
    	    	D2UV:  out Vec from gp);
		     
    	---Purpose: Returns all first and second derivatives.
    
    

    Tolerance(myclass; Quad: Quadric from IntSurf )
    
	---Purpose: returns the tolerance of the zero of the implicit function

    	returns Real from Standard; 


end QuadricTool;


