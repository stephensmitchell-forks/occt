-- Created on: 1991-09-06
-- Created by: NW,JPB,CAL
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Group from Graphic3d inherits TShared
    
        ---Version:

        ---Purpose: This class allows the definition of groups
        --     of primitives inside of graphic objects (presentations).
        --     A group contains the primitives and attributes
        --     for which the range is limited to this group.
        --     The primitives of a group can be globally suppressed.
        --
        --      There are two main group usage models:
        --
        --        1) Non-modifiable, or unbounded, group ('black box'). 
        --           Developers can repeat a sequence of 
        --           SetPrimitivesAspect() with AddPrimitiveArray() methods arbitrary number of times
        --           to define arbitrary number of primitive "blocks" each having individual apect values.
        --           Any modification of such a group is forbidden, as aspects and primitives are mixed 
        --           in memory without any high-level logical structure, and any modification is very likely to result
        --           in corruption of the group internal data.
        --           It is necessary to recreate such a group as a whole when some attribute should be changed.
        --           (for example, in terms of AIS it is necessary to re-Compute() the whole presentation each time).
        --        2) Bounded group. Developers should specify the necessary group aspects with help of
        --           SetGroupPrimitivesAspect() and then add primitives to the group.
        --           Such a group have simplified organization in memory (a single block of attributes
        --           followed by a block of primitives) and therefore it can be modified, if it is necessary to
        --           change parameters of some aspect that has already been set, using methods:
        --           IsGroupPrimitivesAspectSet() to detect which aspect was set for primitives;
        --           GroupPrimitivesAspect() to read current aspect values
        --           and SetGroupPrimitivesAspect() to set new values.
        -- 
        --        Developers are strongly recommended to take all the above into account when filling Graphic3d_Group
        --        with aspects and primitives and choose the group usage model beforehand out of application needs.

        ---Warning:
        ---References:
    
    uses
    
        Array1OfInteger             from TColStd,
        Array1OfReal                from TColStd,
        HArray1OfByte               from TColStd,
    
        ExtendedString              from TCollection,
    
        PlaneAngle                  from Quantity,

    	GroupAspect	            from Graphic3d,
        AspectLine3d                from Graphic3d,
        AspectMarker3d              from Graphic3d,
        AspectText3d                from Graphic3d,
        AspectFillArea3d            from Graphic3d,
        CAspectLine                 from Graphic3d,
        CAspectFillArea             from Graphic3d,
        CAspectMarker               from Graphic3d,
        CAspectText                 from Graphic3d,
        CStructurePtr               from Graphic3d,
        HorizontalTextAlignment     from Graphic3d,
        CBitFields4                 from Graphic3d,
        GraphicDriver               from Graphic3d,
        Structure                   from Graphic3d,
        StructurePtr                from Graphic3d,
        TextPath                    from Graphic3d,
        Vector                      from Graphic3d,
        Array1OfVertex              from Graphic3d,
        Array2OfVertex              from Graphic3d,
        Vertex                      from Graphic3d,
        VerticalTextAlignment       from Graphic3d,
        ArrayOfPrimitives           from Graphic3d,
        TypeOfPrimitiveArray        from Graphic3d,
        IndexBuffer                 from Graphic3d,
        Buffer                      from Graphic3d,
        BoundBuffer                 from Graphic3d,
        TransModeFlags              from Graphic3d,
        BndBox4f                    from Graphic3d,
        Volume                      from Graphic3d,
        Ax2                         from gp
    
    raises

        GroupDefinitionError        from Graphic3d,

    OutOfRange          from Standard
    
    is
        Initialize (theStructure : Structure from Graphic3d)
            returns Group from Graphic3d;
        ---Level: Public
        ---Purpose: Creates a group in the structure <AStructure>.
    
        ---------------------------------------------------
        -- Category: Methods to modify the class definition
        ---------------------------------------------------
    
        Clear ( me  : mutable;
                theUpdateStructureMgr : Boolean from Standard = Standard_True )
        is virtual;
        ---Level: Public
        ---Purpose: Supress all primitives and attributes of <me>.
        --          To clear group without update in Graphic3d_StructureManager
        --          pass Standard_False as <theUpdateStructureMgr>. This
        --          used on context and viewer destruction, when the pointer
        --          to structure manager in Graphic3d_Structure could be 
        --          already released (pointers are used here to avoid handle 
        --          cross-reference);
        ---Category: Methods to modify the class definition

        UpdateAspectLine ( me          : mutable;
                           theIsGlobal : Boolean from Standard )
        is deferred;

        UpdateAspectFace ( me          : mutable;
                           theIsGlobal : Boolean from Standard )
        is deferred;

        UpdateAspectMarker ( me          : mutable;
                             theIsGlobal : Boolean from Standard )
        is deferred;

        UpdateAspectText ( me          : mutable;
                           theIsGlobal : Boolean from Standard )
        is deferred;

        Destroy ( me    : mutable )
            is static;
        ---Level: Public
        ---Purpose: Supress the group <me> in the structure.
        ---Category: Methods to modify the class definition
        ---C++: alias ~
    
        Remove ( me : mutable )
            is static;
        ---Level: Public
        ---Purpose: Supress the group <me> in the structure.
        --  Warning: No more graphic operations in <me> after this call.
        ---Category: Methods to modify the class definition

        --SetTransformPersistence( me     : mutable;
        --                         AFlag  : TransModeFlags from Graphic3d )
        ---Level: Public
    ---Purpose: Modifies the current modelling transform persistence (pan, zoom or rotate)
        --is static;

    --TransformPersistence( me )
    --      returns TransModeFlags from Graphic3d
        ---Level: Public
    ---Purpose: Get the current modelling transform persistence (pan, zoom or rotate)
        --is static;
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectLine3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the line primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectFillArea3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the face primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectText3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the text primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetGroupPrimitivesAspect ( me   : mutable;
                                   CTX  : AspectMarker3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the context for all the marker primitives
        --      of the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectLine3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the line primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectFillArea3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the face primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectText3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the text primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetPrimitivesAspect ( me    : mutable;
                              CTX   : AspectMarker3d from Graphic3d )
            is static;
        ---Level: Public
        ---Purpose: Modifies the current context of the group to give
        --      another aspect for all the marker primitives created
        --      after this call in the group.
        ---Category: Methods to modify the class definition
    
        SetMinMaxValues ( me                : mutable;
                          XMin, YMin, ZMin  : Real from Standard;
                          XMax, YMax, ZMax  : Real from Standard )
            is static;
        ---Level: Public
        ---Purpose: Sets the coordinates of the boundary box of the
        --      group <me>.
        ---Category: Methods to modify the class definition

        -----------------------------------
        -- Category: Methods to create Text
        -----------------------------------
    
        --------------------------------------------
        -- Summary of Texts                       --
        --                                        --
        -- Text  has  geometric  and nongeometric --
        -- attributes.                            --
        --                                        --
        -- The geometric text attributes are :    --
        --                                        --
        --  Character Height.                 --
        --  Character Up Vector.              --
        --  Text Path.                        --
        --  Text Alignment Horizontal.        --
        --  Text Alignment Vertical.          --
        --                                        --
        -- The nongeometric text attributes are : --
        --                                        --
        --  Text Font.                        --
        --  Character Spacing.                --
        --  Character Expansion Factor.       --
        --  Text Color.                       --
        --------------------------------------------
    
        Text (  me  : mutable;
            AText   : CString from Standard;
            APoint  : Vertex from Graphic3d;
            AHeight : Real from Standard;
            AAngle  : PlaneAngle from Quantity;
            ATp : TextPath from Graphic3d;
            AHta    : HorizontalTextAlignment from Graphic3d;
            AVta    : VerticalTextAlignment from Graphic3d;
            EvalMinMax  : Boolean from Standard = Standard_True )
        is virtual;
        ---Level: Public
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      AAngle  : Orientation of the text
        --            (with respect to the horizontal).
        ---Category: Methods to create Text

        Text ( me   : mutable;
               AText    : CString from Standard;
               APoint   : Vertex from Graphic3d;
               AHeight  : Real from Standard;
               EvalMinMax   : Boolean from Standard = Standard_True )
            is static;
        ---Level: Public
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      The other attributes have the following default values:
        --      AAngle  : PI / 2.
        --      ATp     : TP_RIGHT
        --      AHta    : HTA_LEFT
        --      AVta    : VTA_BOTTOM
        ---Category: Methods to create Text
    
        Text (  me          : mutable;
                AText       : ExtendedString from TCollection;
                APoint      : Vertex from Graphic3d;
                AHeight     : Real from Standard;
                AAngle      : PlaneAngle from Quantity;
                ATp         : TextPath from Graphic3d;
                AHta        : HorizontalTextAlignment from Graphic3d;
                AVta        : VerticalTextAlignment from Graphic3d;
                EvalMinMax  : Boolean from Standard = Standard_True )
            is static;
        ---Level: Internal
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      AAngle  : Orientation of the text
        --            (with respect to the horizontal).
        ---Category: Methods to create Text
    
        Text ( me           : mutable;
               AText        : ExtendedString from TCollection;
               APoint       : Vertex from Graphic3d;
               AHeight      : Real from Standard;
               EvalMinMax   : Boolean from Standard = Standard_True )
            is static;
        ---Level: Internal
        ---Purpose: Creates the string <AText> at position <APoint>.
        --      The 3D point of attachment is projected. The text is
        --      written in the plane of projection.
        --      The attributes are given with respect to the plane of
        --      projection.
        --      AHeight : Height of text.
        --            (Relative to the Normalized Projection
        --              Coordinates (NPC) Space).
        --      The other attributes have the following default values:
        --      AAngle  : PI / 2.
        --      ATp     : TP_RIGHT
        --      AHta    : HTA_LEFT
        --      AVta    : VTA_BOTTOM
        ---Category: Methods to create Text
    
        ---------------------------------------
        ---Category: Methods to create Triangle
        ---------------------------------------

    AddPrimitiveArray (me              : mutable;
                       theType         : TypeOfPrimitiveArray from Graphic3d;
                       theIndices      : IndexBuffer          from Graphic3d;
                       theAttribs      : Buffer               from Graphic3d;
                       theBounds       : BoundBuffer          from Graphic3d;
                       theToEvalMinMax : Boolean from Standard = Standard_True) is virtual;
    ---Level: Public
    ---Purpose: Adds an array of primitives for display

    AddPrimitiveArray( me      : mutable;
                       thePrim : ArrayOfPrimitives from Graphic3d;
                       theToEvalMinMax : Boolean from Standard = Standard_True );
    ---Level: Public
    ---Purpose: Adds an array of primitives for display

    AddVolume (me              : mutable;
               theVolume       : Volume from Graphic3d;
               theToEvalMinMax : Boolean from Standard = Standard_True) is virtual;
    ---Level: Public
    ---Purpose: Adds volume of voxels for display

    Marker ( me              : mutable;
             thePoint        : Vertex from Graphic3d;
             theToEvalMinMax : Boolean from Standard = Standard_True )
    is static;
    ---Level: Public
    ---Purpose: Creates a primitive array with single marker using AddPrimitiveArray().

    UserDraw ( me               : mutable;
               theObject        : Address from Standard;
               theToEvalMinMax  : Boolean from Standard = Standard_True;
               theContainsFacet : Boolean from Standard = Standard_False )
    is virtual;
    ---Level: Public
    ---Purpose: Creates a UserDraw primitive using obsolete API.

    SetStencilTestOptions (me          : mutable;
                           theIsEnabled: Boolean from Standard)
    is deferred;
    ---Purpose: sets the stencil test to theIsEnabled state;

    SetFlippingOptions (me           : mutable;
                        theIsEnabled : Boolean from Standard;
                        theRefPlane  : Ax2 from gp)
    is deferred;
    ---Purpose: sets the flipping to theIsEnabled state.

        ----------------------------
        -- Category: Inquire methods
        ----------------------------

        IsGroupPrimitivesAspectSet ( me;
                    theAspect : GroupAspect from Graphic3d )
            returns Boolean from Standard
            is static;
        ---Level: Public
        ---Purpose: Returns TRUE if aspect is set for the group.
        ---Category: Inquire methods

    	GroupPrimitivesAspect ( me;
    				CTXL	: AspectLine3d from Graphic3d;
    				CTXT	: AspectText3d from Graphic3d;
    				CTXM	: AspectMarker3d from Graphic3d;
    				CTXF	: AspectFillArea3d from Graphic3d )
    		is static;
    	---Level: Public
    	---Purpose: Returns the context of all the primitives of the group.
    	---Category: Inquire methods
    
    	PrimitivesAspect ( me;
    			   CTXL	: AspectLine3d from Graphic3d;
    			   CTXT	: AspectText3d from Graphic3d;
    			   CTXM	: AspectMarker3d from Graphic3d;
    			   CTXF	: AspectFillArea3d from Graphic3d )
    		is static;
    	---Level: Public
    	---Purpose: Returns the last inserted context in the group <me>
    	--	    foreach kind of primitives.
    	---Category: Inquire methods

        ContainsFacet ( me )
            returns Boolean from Standard
            is static;
        ---Level: Internal
        ---Purpose: Returns Standard_True if the group <me> contains
        --      Polygons, Triangles or Quadrangles.
        ---Category: Inquire methods
    
        IsDeleted ( me )
            returns Boolean from Standard
            is static;
        ---Level: Public
        ---Purpose: Returns Standard_True if the group <me> is deleted.
        --      <me> is deleted after the call Remove (me) or the
        --      associated structure is deleted.
        ---Category: Inquire methods
    
        IsEmpty ( me )
            returns Boolean from Standard
            is static;
        ---Level: Public
        ---Purpose: Returns Standard_True if the group <me> is empty.
        ---Warning: A group is empty if the MinMaxValues method returns :
        --      XMin = YMin = ZMin = RealFirst ().
        --      XMax = YMax = ZMax = RealLast ().
        ---Category: Inquire methods
    
        MinMaxValues ( me;
                       XMin, YMin, ZMin : out Real from Standard;
                       XMax, YMax, ZMax : out Real from Standard )
            is static;
        ---Level: Public
        ---Purpose: Returns the coordinates of the boundary box of the
        --      group <me>.
        ---Warning: If the group <me> is empty then :
        --      XMin = YMin = ZMin = RealFirst ().
        --      XMax = YMax = ZMax = RealLast ().
        ---Category: Inquire methods

        BoundingBox ( me )
            returns BndBox4f from Graphic3d
            is static;
        ---Level: Public
        ---Purpose: Returns boundary box of the group <me> without transformation applied,
        ---if it is specified for the structure.
        ---C++: return const &

        ChangeBoundingBox ( me : mutable )
            returns BndBox4f from Graphic3d
            is static;
        ---Level: Public
        ---Purpose: Returns non-const boundary box of the group <me> without transformation applied,
        ---if it is specified for the structure.
        ---C++: return &
    
        Structure ( me )
            returns Structure from Graphic3d
            is static;
        ---Level: Public
        ---Purpose: Returns the structure containing the group <me>.
        ---Category: Inquire methods
    
        ----------------------------
        -- Category: Private methods
        ----------------------------
        
        MinMaxCoord ( me;
                      XMin, YMin, ZMin : out Real from Standard;
                      XMax, YMax, ZMax : out Real from Standard )
            is static private;
        ---Level: Internal
        ---Purpose: Returns the extreme coordinates found in the group.
        ---Warning: If the group <me> is empty then :
        --      XMin = YMin = ZMin = RealFirst ().
        --      XMax = YMax = ZMax = RealLast ().
        ---Category: Private methods
    
        Update ( me )
            is static private;
        ---Level: Internal
        ---Purpose: Calls the Update method of the StructureManager which
        --      contains the associated Structure of the Group <me>.
        ---Category: Private methods

        SetClosed (me: mutable; theIsClosed : Boolean from Standard);
        ---Purpose: Changes property shown that primitive arrays within this group form closed volume (do no contain open shells).

        IsClosed (me) returns Boolean from Standard;
        ---Purpose: Return true if primitive arrays within this graphic group form closed volume (do no contain open shells).

    fields
    
    --
    -- Class    :   Graphic3d_Group
    --
    -- Purpose  :   Declaration of variables specific to groups
    --          of primitives.
    --
    -- Reminder :   A group is defined in a structure
    --          It acts as the smallest editable entity.

  -- the state of the different contexts for primitives
  myCBitFields   : CBitFields4 from Graphic3d is protected;

  -- the structure contains the group
  myStructure    : StructurePtr from Graphic3d is protected;

  -- the min-max
  myBounds        : BndBox4f from Graphic3d is protected;

  -- Identifies group forming closed volume. Used to filter groups for back face culling and capping algorithms.
  myIsClosed  : Boolean from Standard is protected;

  ContextLine     : CAspectLine     from Graphic3d is protected;
  ContextFillArea : CAspectFillArea from Graphic3d is protected;
  ContextMarker   : CAspectMarker   from Graphic3d is protected;
  ContextText     : CAspectText     from Graphic3d is protected;

friends

  class Structure from Graphic3d

end Group;
