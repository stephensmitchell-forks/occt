-- Created on: 1994-11-25
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Builder from TopoDSToStep
    inherits Root from TopoDSToStep

    ---Purpose: This builder Class provides services to build
    --          a ProSTEP Shape model from a Cas.Cad BRep.                 

uses

    FinderProcess_Handle          from Transfer,
    Shape                         from TopoDS,
    Tool                          from TopoDSToStep,
    BuilderError                  from TopoDSToStep,
    TopologicalRepresentationItem from StepShape

raises NotDone from StdFail 
    
is 

--  -----------------------------------------------------------
--  Constructor
--  -----------------------------------------------------------

    Create returns Builder from TopoDSToStep;
    
    Create(S           : Shape from TopoDS;
           T           : in out Tool from TopoDSToStep;
           FP          : FinderProcess_Handle from Transfer)
    	returns Builder from TopoDSToStep;
    
    Init(me          : in out;
         S           : Shape from TopoDS;
         T           : in out Tool from TopoDSToStep;
         FP          : FinderProcess_Handle from Transfer);
    
--  -----------------------------------------------------------    
--  Get the Result
--  -----------------------------------------------------------

    Error(me) returns BuilderError from TopoDSToStep;
    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const &

fields

    myResult : TopologicalRepresentationItem from StepShape;
    
    myError  : BuilderError                  from TopoDSToStep;

end Builder;
