-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentRetrievalDriver from XmlLDrivers inherits RetrievalDriver from PCDM

uses
    ExtendedString		from TCollection,
    SequenceOfExtendedString	from TColStd,
    Document			from PCDM,
    Document			from CDM,
    Document			from TDocStd,
    IODevice          from Storage,
    Application			from CDM,
    ADriver		        from XmlMDF, 
    ADriverTable		from XmlMDF,
    RRelocationTable		from XmlObjMgt,
    Element			from XmlObjMgt,
    MessageDriver               from CDM

is
    Create returns DocumentRetrievalDriver from XmlLDrivers;
    -- Constructor

    SchemaName		(me)
	returns ExtendedString from TCollection is redefined virtual;
    -- pure virtual method definition

    Make		(me : mutable; PD : Document from PCDM;
				       TD : Document from CDM)
	is redefined virtual;
    -- pure virtual method definition

    CreateDocument	(me : mutable)
	returns Document from CDM is redefined virtual;
    -- pure virtual method definition

    Read(me:mutable; theDevice: IODevice from Storage;
    	    	     theNewDocument: Document    from CDM;
    	    	     theApplication: Application from CDM) is redefined virtual;
    -- 

    ReadFromDomDocument (me : mutable; theDomElement: Element from XmlObjMgt;
				       theNewDocument: Document from CDM;
				       theApplication: Application from CDM)
	is virtual protected;

    MakeDocument	(me : mutable; thePDoc: Element  from XmlObjMgt;
    	    	    	       theTDoc: Document from CDM)
    	returns Boolean from Standard
	is virtual protected;

    AttributeDrivers	(me : mutable; theMsgDriver: MessageDriver from CDM)
	returns ADriverTable from XmlMDF
	is virtual; 
	
    ReadShapeSection (me:mutable; thePDoc  :  Element from XmlObjMgt; 
    	    	    	    	  theMsgDriver : MessageDriver from CDM) 
        returns ADriver from XmlMDF
        is virtual protected; 
	 
    ShapeSetCleaning(me:mutable; theDriver : ADriver from XmlMDF) 
        is virtual protected;  
	
    PropagateDocumentVersion(me:mutable; theDocVersion : Integer from Standard) 
        is virtual protected; 
	
fields
    myDrivers	: ADriverTable		from XmlMDF      is protected;
    myRelocTable: RRelocationTable	from XmlObjMgt   is protected;
    myDevice  : IODevice from Storage is protected;

end DocumentRetrievalDriver;
