-- Created on: 1994-11-25
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package TopoDSToStep

    ---Purpose: This package implements the mapping between CAS.CAD
    --  Shape representation and AP214 Shape Representation.
    --  The target schema is pms_c4 (a subset of AP214)
    --  
    --  How to use this Package :
    --  
    --  Entry point are context dependent. It can be :
    --     MakeManifoldSolidBrep
    --     MakeBrepWithVoids
    --     MakeFacetedBrep
    --     MakeFacetedBrepAndBrepWithVoids
    --     MakeShellBasedSurfaceModel
    --  Each of these classes call the Builder
    --  The class tool centralizes some common informations.   

uses TopoDS, StdFail, TCollection, TColStd, TopTools, Transfer, MoniTool,
     BRepTools, TopLoc, GeomAbs, Geom2d, Geom, gp,
     StepGeom, StepShape

is

--  ------------------------------------------------------
--  Enumeration
--  ------------------------------------------------------

    enumeration BuilderError is
    	BuilderDone,
	NoFaceMapped,
	BuilderOther
    end BuilderError;
    
    enumeration MakeFaceError is
    	FaceDone,
	InfiniteFace,
	NonManifoldFace,
	NoWireMapped,
    	FaceOther
    end MakeFaceError;
    
    enumeration MakeWireError is
    	WireDone,
	NonManifoldWire,
    	WireOther
    end MakeWireError;
    
    enumeration MakeEdgeError is
    	EdgeDone,
	NonManifoldEdge,
    	EdgeOther
    end MakeEdgeError;
    
    enumeration MakeVertexError is
    	VertexDone,
    	VertexOther
    end MakeVertexError;
    
    enumeration FacetedError is
	FacetedDone,    
    	SurfaceNotPlane,
	PCurveNotLinear
    end FacetedError;

--  ------------------------------------------------------
--  Package Classes
--  ------------------------------------------------------

    private deferred class Root;

    class MakeManifoldSolidBrep;

    class MakeBrepWithVoids;

    class MakeFacetedBrep;

    class MakeFacetedBrepAndBrepWithVoids;

    class MakeShellBasedSurfaceModel;

    class MakeGeometricCurveSet;
    
    class Builder;
    
    class WireframeBuilder;
    
    class Tool;
    
    class FacetedTool;
    
    class MakeStepFace;
    
    class MakeStepWire;
    
    class MakeStepEdge;
    
    class MakeStepVertex;
    
--    private class DirectModification;
--    private class ConicalSurfModif;
    
--  ------------------------------------------------------
--  Instanciated Class
--  ------------------------------------------------------

--    class DataMapOfShape instantiates
--    	  DataMap from TCollection 
--    	    (Shape                         from TopoDS,
--    	     TopologicalRepresentationItem from StepShape,
--	     ShapeMapHasher                from TopTools);

--  ------------------------------------------------------
--  Package Method
--  ------------------------------------------------------

    DecodeBuilderError(E : BuilderError from TopoDSToStep)
    	returns HAsciiString from TCollection;   
   
    DecodeFaceError(E : MakeFaceError from TopoDSToStep)
    	returns HAsciiString from TCollection;
	
    DecodeWireError(E : MakeWireError from TopoDSToStep)
    	returns HAsciiString from TCollection;   
   
    DecodeEdgeError(E : MakeEdgeError from TopoDSToStep)
    	returns HAsciiString from TCollection;
	
    DecodeVertexError(E : MakeVertexError from TopoDSToStep)
    	returns HAsciiString from TCollection;
	
--    DirectFaces(S : Shape from TopoDS)
--    	returns Shape from TopoDS;
	---Purpose: Returns a new shape without undirect surfaces.
	
    AddResult (FP: FinderProcess_Handle from Transfer;
     	       Shape: Shape from TopoDS;
	       entity: Transient from Standard);
	---Purpose: Adds an entity into the list of results (binders) for
	--          shape stored in FinderProcess

    AddResult (FP: FinderProcess_Handle from Transfer;
     	       Tool: Tool from TopoDSToStep);
	---Purpose: Adds all entities recorded in Tool into the map of results
	--          (binders) stored in FinderProcess

end TopoDSToStep;
