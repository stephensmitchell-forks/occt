-- File:	Unfolding.cdl
-- Created:	Tue Jul 22 12:48:05 2008
-- Author:	Sergey KHROMOV
--		<skv@dimox>
---Copyright:	Open CASCADE 2008

package Unfolding
    ---Purpose: This package contains a tool for unfolding a surface on a plane.

uses

    TopoDS,
    TopTools,
    gp,
    Standard,
    TCollection,
    TColgp,
    math

is

    ---Purpose: Enumeration that defines an error status of an operation.
    enumeration ErrorStatus
    is
    	Done,
	NotDone,
	Failure,
	InvalidSurface,
	InvalidInput,
	InvalidShape,
	ComplexShape
    end;

    class Surface;

    class Point;
    
    class FunctionWithDerivative;
    
    class Shell;

    class FaceDataContainer;

    class FaceDataMapHasher;

    class Array2OfPoint
          instantiates Array2 from TCollection (Point from Unfolding);

    class HArray2OfPoint
    	instantiates HArray2 from TCollection (Point         from Unfolding,
    	    	    	    	    	       Array2OfPoint from Unfolding);

    class IndexedMapOfFaceDataContainer
    	instantiates IndexedMap from TCollection
                                           (FaceDataContainer from Unfolding,
                                            FaceDataMapHasher from Unfolding);

    ToShell(theShape     :     Shape       from TopoDS;
            theTolerance :     Real        from Standard;
            theStatus    : out ErrorStatus from Unfolding)
    ---Purpose: This method converts theShape to a shell. It sewes faces of the
    --          shell if it is necessary and possible with the given tolerance.
    --          If it is not possible to construct a single shell from theShape,
    --          this method returns null shell and the corresponding error
    --          status. The status can have the following values:
    --            -  Unfolding_Done: the operation succeeded
    --            -  Unfolding_InvalidInput: input shape type is less then
    --                  TopAbs_SHELL.
    --            -  Unfolding_Failure: sewing failure.
    --            -  Unfolding_InvalidShape: the shape after sewing does not
    --                   contain shells.
    --            -  Unfolding_ComplexShape: the shape after sewing contains
    --                   either more then one shell or one shell and other not
    --                   connected shapes.
    returns Shell from TopoDS;

    NbSamples(theEdge     : Edge        from TopoDS;
    	      theFaces    : ListOfShape from TopTools;
    	      theTolerance: Real        from Standard)
    ---Purpose: This method returns the number of sample points for theEdge.
    --          theFaces is a list of faces that contain theEdge.
    returns Integer from Standard;

    GetMaxNbSamples
    ---Purpose: This method returns the maximal number of points for sampling of
    --          edges and/or faces.
    ---C++: inline
    returns Integer from Standard;

end Unfolding;
