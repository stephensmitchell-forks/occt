-- Created on: 2000-09-28
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ExternFile from STEPCAFControl inherits TShared from MMgt

    ---Purpose: Auxiliary class serving as container for data resulting
    --          from translation of external file

uses
    HAsciiString from TCollection,
    ReturnStatus from IFSelect,
    WorkSession_Handle from XSControl,
    Shape from TopoDS,
    Label from TDF

is

    Create returns ExternFile;
    	---Purpose: Creates an empty structure
	
    SetWS (me: mutable; WS: WorkSession_Handle from XSControl);
    	---C++: inline
    GetWS (me) returns WorkSession_Handle from XSControl;
    	---C++: inline
    
    SetLoadStatus (me: mutable; stat: ReturnStatus from IFSelect);
    	---C++: inline
    GetLoadStatus (me) returns ReturnStatus from IFSelect;
    	---C++: inline
    
    SetTransferStatus (me: mutable; isok: Boolean);
    	---C++: inline
    GetTransferStatus (me) returns Boolean;
    	---C++: inline
    
    SetWriteStatus (me: mutable; stat: ReturnStatus from IFSelect);
    	---C++: inline
    GetWriteStatus (me) returns ReturnStatus from IFSelect;
    	---C++: inline
    
    SetName (me: mutable; name: HAsciiString from TCollection);
    	---C++: inline
    GetName (me) returns HAsciiString from TCollection;
    	---C++: inline
    
--    SetShape (me: mutable; S: Shape from TopoDS);
    	---C++: inline
--    GetShape (me) returns Shape from TopoDS;
    	---C++: inline
    
    SetLabel (me: mutable; L: Label from TDF);
    	---C++: inline
    GetLabel (me) returns Label from TDF;
    	---C++: inline
    
fields

    myWS   : WorkSession_Handle from XSControl;
    
    myLoadStatus: ReturnStatus from IFSelect;
    myTransferStatus: Boolean;
    myWriteStatus: ReturnStatus from IFSelect;

    myName: HAsciiString from TCollection;

--    myShape: Shape from TopoDS;
    myLabel: Label from TDF;

end ExternFile;
