-- Created by: Peter KURNEV
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BOPAlgo 
---Purpose: 

uses
    gp,  
    Bnd, 
    Message,
    TopAbs, 
    Geom,  
    GeomAPI, 
    BRepClass3d,
    TopoDS, 
    TopTools, 
    IntTools,
    IntSurf,
    --
    BOPDS, 
    BOPCol, 
    BOPTools 
is   
    enumeration Operation is  
      COMMON, 
      FUSE, 
      CUT,    
      CUT21,
      SECTION, 
      UNKNOWN
    end Operation;   
     
    enumeration CheckStatus is
      CheckUnknown,
      BadType,
      SelfIntersect,
      TooSmallEdge,
      NonRecoverableFace,
      IncompatibilityOfVertex,
      IncompatibilityOfEdge,
      IncompatibilityOfFace, 
      OperationAborted,
      GeomAbs_C0,
      InvalidCurveOnSurface,
      NotValid
    end CheckStatus;

    --
    -- classes 
    --   
    deferred class Algo; 
    deferred class BuilderShape; 
    class PaveFiller;
    class Builder; 
    class BOP;   
    class Section;   
    --	
    deferred class BuilderArea;
    class BuilderFace;
    class WireEdgeSet;
    class WireSplitter;  
    class ShellSplitter;  
    class BuilderSolid; 
    class Tools; 
    class SectionAttribute; 
    class CheckerSI; 
    class ArgumentAnalyzer; 
    class CheckResult; 
    class MakerVolume;
    --
    --  pointers
    --
    pointer PPaveFiller to PaveFiller from BOPAlgo; 
    pointer PWireEdgeSet to WireEdgeSet from BOPAlgo;  
    pointer PSection to Section from BOPAlgo;   
    pointer PBOP to BOP from BOPAlgo;  
    pointer PBuilder to Builder from BOPAlgo;  
    pointer PArgumentAnalyzer to ArgumentAnalyzer from BOPAlgo;  
    -- 
    imported ListOfCheckResult; 
    imported CellsBuilder;
    
end BOPAlgo;
