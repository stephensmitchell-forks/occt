-- Created on: 1997-08-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Application from CDF inherits Application from CDM

uses  
    ExtendedString from TCollection,  
    ExtendedString from TCollection,  
    Document from CDM,  
    Manager from Resource, 
    MetaData from CDM,  
    ReaderStatus  from PCDM,  
    GUID from Standard, 
    Reader from PCDM,  
    Writer from PCDM, 
    TypeOfActivation from CDF, 
    SequenceOfExtendedString from TColStd, 
    CanCloseStatus from CDM,  
    AsciiString from TCollection,
    IODevice from Storage
    
raises NoSuchObject from Standard
is


    Initialize;
    
    Load(myclass; aGUID:GUID from Standard)
    returns  mutable Application from CDF;
    ---Purpose: plugs an application.
    

---Category: Open closing of documents
---Purpose:
-- Open is used 
--       - for opening a Document that has been created in an application
--       - for opening a Document from the database
--       - for opening a Document from a file.
--  The Open methods always add the document in the session directory and 
--  calls the virtual Activate method. The document is considered to be 
--  opened until Close is used. To be storable, a document must be 
--  opened by an application since the application resources are 
--  needed to store it.
--          
--          
--          
--          
    Open(me: mutable; aDocument: Document from CDM);
    ---Purpose: puts the document in the current session directory
    --          and calls the virtual method Activate on it.
    
    
    CanClose(me: mutable; aDocument: Document from CDM)
    returns CanCloseStatus from CDM;
    
    Close(me: mutable; aDocument: Document from CDM);
    ---Purpose: removes the document of the current session directory 
    --          and closes the document;
    
    Retrieve (me: mutable; aDevice: in out IODevice from Storage; UseStorageConfiguration: Boolean from Standard = Standard_True)
    returns Document from CDM;
    ---Purpose: This method retrieves a document from the database. 
    --          If the Document references other documents which have
    --          been updated, the latest version of these documents will 
    --          be used if {UseStorageConfiguration} is Standard_True.
   --           The content of {aFolder}, {aName} and {aVersion} depends on 
   --           the Database Manager system. If the DBMS is only based on 
   --           the OS, {aFolder} is a directory and {aName} is the name of a 
   --           file. In this case the use of the syntax with {aVersion} 
   --           has no sense. For example: 
--
-- Handle(CDM_Document) theDocument=myApplication->Retrieve("/home/cascade","box.dsg");
--              If the DBMS is EUCLID/Design Manager, {aFolder}, {aName} 
--              have the form they have in EUCLID/Design Manager. For example:
--              
-- Handle(CDM_Document) theDocument=myApplication->Retrieve("|user|cascade","box"); 
-- 
-- Since  the version is not specified in  this syntax, the  latest wil be used.
--  A link is kept with the database through an instance of CDM_MetaData


    Retrieve (me: mutable; aDevice: in out IODevice from Storage; aVersion: ExtendedString from TCollection; UseStorageConfiguration: Boolean from Standard = Standard_True)
    returns Document from CDM;
    ---Purpose:  This method retrieves  a  document from the database.
    --          If the  Document references other documents which have
    --          been  updated, the  latest version of  these documents
    --           will    be   used  if   {UseStorageConfiguration}  is
    --          Standard_True.  --  If the DBMS is  only  based on the
    --           OS, this syntax  should not be used.
    --           
--              If the DBMS is EUCLID/Design Manager, {aFolder}, {aName} 
--              and  {aVersion} have the form they have in 
--              EUCLID/Design Manager. For example:
--              
-- Handle(CDM_Document) theDocument=myApplication->Retrieve("|user|cascade","box","2");
--             A link is kept with the database through an instance 
--             of CDM_MetaData

    CanRetrieve(me: mutable; aDevice: in out IODevice from Storage)
    ---Purpose:
    returns ReaderStatus from PCDM;
    
    CanRetrieve(me: mutable; aDevice: in out IODevice from Storage; aVersion: ExtendedString from TCollection)
    ---Purpose:
    returns ReaderStatus from PCDM;

    Formats(me: mutable; Formats: out SequenceOfExtendedString from TColStd) 
    is deferred;

---Category: CurrentDocument methods.
--           

    GetRetrieveStatus(me) returns ReaderStatus from PCDM; 
    ---C++: inline     
    ---Purpose: Checks  status  after  Retrieve 
     
   ---Category: Store&Retrieve virtuals methods

    Activate(me: mutable; aDocument: Document from CDM; aTypeOfActivation: TypeOfActivation from CDF)
    is virtual private;
    ---Purpose: Informs the  application that aDocument has  been
    --          activated. A document is activated when it is created or 
    --          retrieved.
    --    aTypeOfActivation will be:
    --            - CDF_TOA_New if the document is a new one 
    --              (even empty or retrieved from the database for 
    --              the first time).
    --            - CDF_TOA_Unchanged if the document was already 
    --              retrieved but had no changes since the previous retrieval.
    --            - CDF_TOA_Modified if the document was already 
    --              retrieved and modified since the previous retrieval.
    --  You do not need to call <Activate>, but you should  redefine 
    --  this method to implement application specific behavior.


 ---Category:  methods to get storage/retrieval driver.
 --           
 --           
    FindReader(me: mutable; aDevice: IODevice from Storage)
    returns Boolean from Standard;

    Reader(me: mutable; aDevice: IODevice from Storage) 
    returns Reader from PCDM
    raises NoSuchObject from Standard;
    
    FindReaderFromFormat(me: mutable; aFormat: ExtendedString from TCollection)
    returns Boolean from Standard;
    
    ReaderFromFormat(me: mutable; aFormat: ExtendedString from TCollection) 
    returns Reader from PCDM
    raises NoSuchObject from Standard;

    ---Purpose: 

    Format (me : mutable; aDevice : IODevice from Storage; 
                          theFormat : out ExtendedString from TCollection)
    ---Purpose: try to  retrieve a Format  directly in the  file or in
    --           application   resource  by using   extension. returns
    --          True if found;
    returns Boolean from Standard;
    
---Category: Default Storage folder
--           
    DefaultFolder(me: mutable) returns ExtString from Standard;
    
    SetDefaultFolder(me: mutable; aFolder: ExtString from Standard)
    returns Boolean from Standard;
    
    DefaultExtension(me: mutable) returns ExtString from Standard;
    
---Category: private methods
    Retrieve(me: mutable; aMetaData: MetaData from CDM; UseStorageConfiguration: Boolean from Standard)
    returns mutable Document from CDM
    is private;

    Retrieve(me: mutable; aMetaData: MetaData from CDM; UseStorageConfiguration: Boolean from Standard; IsComponent: Boolean from Standard)
    returns mutable Document from CDM
    is private;

    DocumentVersion(me: mutable; theMetaData: MetaData from CDM)
    returns Integer from Standard
    is private;

    FindReader(me: mutable; aDevice: IODevice from Storage; PluginIn: out GUID from Standard; ResourceName: out ExtendedString from TCollection)
    returns Boolean from Standard
    is private;
    

    FindReaderFromFormat(me: mutable; aFormat: ExtendedString from TCollection; PluginIn: out GUID from Standard; ResourceName: out ExtendedString from TCollection)
    returns Boolean from Standard
    is private;
    
    TypeOfActivation(me: mutable; aMetaData: MetaData from CDM)
    returns TypeOfActivation from CDF
    is private;

    CanRetrieve(me: mutable; aMetaData: MetaData from CDM)
    returns ReaderStatus from PCDM
    is private;
    
fields

    myDefaultFolder: ExtendedString from TCollection; 
    myRetrievableStatus :  ReaderStatus from PCDM  is protected; 
    
friends 
    class Session from CDF--,
    --class CheckDocumentToStore from CDF 

end Application from CDF;
