-- Created on: 1998-09-30
-- Created by: Denis PASCAL
-- Copyright (c) 1998-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Presentation from TDataXtd inherits Attribute from TDF

---Purpose: An attribute to associate an
-- AIS_InteractiveObject to a label in an AIS viewer.
-- This attribute works in collaboration with TPrsStd_AISViewer.
-- Note that all the Set... and Unset... attribute
-- methods as well as the query methods for
-- visualization attributes and the HasOwn... test
-- methods are shortcuts to the respective
-- AIS_InteractiveObject settings.

uses GUID                 from Standard,
     AttributeIndexedMap  from TDF,
     DataSet              from TDF,
     AttributeDelta       from TDF,
     Label                from TDF,
     RelocationTable      from TDF

is

    Create returns Presentation from TDataXtd;
    ---Purpose: Default constructor.

    Set(myclass; theLabel : Label from TDF; theDriverId : GUID from Standard)
    returns Presentation from TDataXtd;
    ---Purpose: Creates or retrieves the presentation attribute on
    -- the label, and sets the GUID driver.

    Set(myclass; theMaster : Attribute from TDF) returns Presentation from TDataXtd;
    ---Purpose:  Creates or retrieves the presentation attribute attached to master.
    -- The GUID of the driver will be the GUID of master.
    -- Master is the attribute you want to display.

    Unset(myclass; theLabel : Label from TDF);
    ---Purpose: Delete (if exist) the presentation attribute associated to the input label.

    GetID(myclass) returns GUID from Standard;
    ---Purpose: Returns the GUID for TDataXtd_Presentation attributes.
    ---C++: return const &

    GetDriverGUID(me) returns GUID from Standard;

    SetDriverGUID(me: mutable ; theGUID : GUID from Standard);

    ID(me)returns GUID from Standard;
    ---C++: return const &


    IsDisplayed(me) returns Boolean from Standard;    
    ---Purpose: Returns true if this presentation attribute is displayed.

    IsHasOwnMaterial(me) returns Boolean from Standard;
    ---Purpose: Returns true if this presentation attribute already has a material setting.

    IsHasOwnTransparency(me) returns Boolean from Standard;
    ---Purpose: Returns true if this presentation attribute already has a transparency setting.

    IsHasOwnColor(me) returns Boolean from Standard;
    ---Purpose: Returns true if this presentation attribute already has a color setting.

    IsHasOwnWidth(me) returns Boolean from Standard;
    ---Purpose: Returns true if this presentation attribute already has a width setting.

    IsHasOwnMode(me) returns Boolean from Standard;

    IsHasOwnSelectionMode(me) returns Boolean from Standard;


    SetDisplayed(me : mutable; theIsDisplayed : Boolean from Standard);

    SetMaterial(me : mutable; theName : Integer from Standard);
    ---Purpose: Sets the material for this presentation  attribute.

    SetTransparency(me : mutable; theValue : Real from Standard = 0.6);
    ---Purpose:
    -- Sets the transparency value for this presentation attribute.
    -- @param theValue - parameter of transparency, this value is 0.6 by default.

    SetColor(me: mutable; theColor : Integer from Standard);
    ---Purpose: Sets the color aColor for this presentation attribute.

    SetWidth(me: mutable; theWidth : Real from Standard);
    ---Purpose: Sets the width for this presentation attribute.

    SetMode(me: mutable; theMode : Integer from Standard);

    SetSelectionMode(me: mutable; theSelectionMode : Integer from Standard);


    Material(me) returns Integer from Standard;
    ---Purpose: Returns the material setting for this presentation attribute.

    Transparency(me) returns Real from Standard;

    Color(me) returns Integer from Standard;

    Width(me) returns Real from Standard;

    Mode(me)  returns  Integer  from  Standard;

    SelectionMode(me) returns Integer from Standard;


    UnsetMaterial(me : mutable);
    ---Purpose: Removes the material setting from this presentation attribute.

    UnsetTransparency(me : mutable);
    ---Purpose: Removes the transparency setting from this presentation attribute.

    UnsetColor(me : mutable);
    ---Purpose: Removes the color setting from this presentation attribute.

    UnsetWidth(me : mutable);
    ---Purpose: Removes the width setting from this presentation attribute.

    UnsetMode(me : mutable);

    UnsetSelectionMode(me : mutable);


    NewEmpty(me) returns Attribute from TDF;

    Restore(me: mutable; theAttribute : Attribute from TDF);

    Paste(me; theInto : Attribute from TDF; theRT : RelocationTable from TDF);

    BackupCopy(me) returns Attribute from TDF is redefined;

fields

    myDriverGUID           : GUID                 from Standard;    
    myColor                : Integer              from Standard;
    myMaterial             : Integer              from Standard;
    myMode                 : Integer              from Standard;
    mySelectionMode        : Integer              from Standard;
    myTransparency         : Real                 from Standard;
    myWidth                : Real                 from Standard;
    myIsDisplayed          : Boolean              from Standard; 
    myIsHasOwnColor        : Boolean              from Standard;
    myIsHasOwnMaterial     : Boolean              from Standard;
    myIsHasOwnTransparency : Boolean              from Standard;    
    myIsHasOwnWidth        : Boolean              from Standard;  
    myIsHasOwnMode         : Boolean              from Standard;
    myIsHasOwnSelectionMode: Boolean              from Standard;

end Presentation;