-- Created on: 1997-08-07
-- Created by: VAUTHIER Jean-Claude 
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- modified     Sergey Zaritchny



package MDataXtd 

	---Purpose: Storage    and  Retrieval  drivers   for modelling
	--          attributes.   Transient  attributes are defined in
	--          package TDataStd and persistent one are defined in
	--          package PDataStd

uses TDF,
     PDF,
     MDF, 
     CDM,
     TDataStd, 
     TDataXtd,
     Geom,  -- a supprimer des que Translate est poussee dans MgtGeom
     PGeom  -- a supprimer des que Translate est poussee dans MgtGeom

is

    	---Purpose: Storage drivers for TDataXtd attributes
    	--          =======================================

        class ShapeStorageDriver;
	
	class PointStorageDriver;
	
	class AxisStorageDriver;
	
	class PlaneStorageDriver;

    	class GeometryStorageDriver;

	class ConstraintStorageDriver;
	
	class PlacementStorageDriver;
	
	class PatternStdStorageDriver;

        class PresentationStorageDriver;

        class PositionStorageDriver;
 
    
    	---Purpose: Retrieval drivers for PDataXtd attributes
    	--          =========================================

	class ShapeRetrievalDriver;	
	
	class PointRetrievalDriver;
	
	class AxisRetrievalDriver;
	
	class PlaneRetrievalDriver;

    	class GeometryRetrievalDriver;

	class ConstraintRetrievalDriver;
	
	class PlacementRetrievalDriver;
	
	class PatternStdRetrievalDriver;

	class PresentationRetrievalDriver;

	class PresentationRetrievalDriver_1;
	
	class PositionRetrievalDriver;



    AddStorageDrivers(aDriverSeq : ASDriverHSequence from MDF; theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute storage drivers to <aDriverSeq>.


    AddRetrievalDrivers(aDriverSeq : ARDriverHSequence from MDF; theMessageDriver : MessageDriver from CDM);
	---Purpose: Adds the attribute retrieval drivers to <aDriverSeq>.


    Translate (Geometry : Geometry from Geom)
    	---Purpose: Method to launch in MgtGeom
    	--           Delete MDataStd_1.cxx
    	--           Modify MDataStd_GeometryStorageDriver::Paste
    returns Geometry from PGeom;


    Translate (Geometry : Geometry from PGeom)
    	---Purpose : Method to lasunch in MgtGeom
    	--           Delete MDataStd_1.cxx
    	--           Modify MDataStd_GeometryRetrievalDriver::Paste
    returns Geometry from Geom;


    ---Purpose: Translation of TDataXtd enumerations to integer
    --          ===============================================
 
    ConstraintTypeToInteger (e : ConstraintEnum from TDataXtd)
    returns Integer from Standard;

    IntegerToConstraintType (i : Integer from Standard)
    returns ConstraintEnum from TDataXtd;     
    
    GeometryTypeToInteger (e : GeometryEnum from TDataXtd)
    returns Integer from Standard;

    IntegerToGeometryType (i : Integer from Standard)
    returns GeometryEnum from TDataXtd;     
    
end MDataXtd;
