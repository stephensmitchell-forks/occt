-- Created on: 1993-10-14
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class BooleanOperation from BRepAlgoAPI
    inherits BuilderAlgo from BRepAlgoAPI
    
    ---Purpose:  
    -- The abstract class BooleanOperation is the root
    -- class of Boolean Operations (see Overview).
    -- Boolean Operations algorithm is divided onto two parts.
    -- - The first one is computing interference between arguments.
    -- - The second one is building the result of operation.
    -- The class BooleanOperation provides API level of both parts
  
uses

    Shape from TopoDS, 
    DataMapOfShapeShape from TopTools, 
    ListOfShape from TopTools, 
    ListOfShape from BOPCol,    
    --
    Operation   from BOPAlgo,
    PaveFiller from BOPAlgo 
    
    
is 
    Initialize
        returns BooleanOperation from BRepAlgoAPI; 
    ---Purpose:  Empty constructor        
     
    Initialize (PF :PaveFiller from BOPAlgo) 
        returns BooleanOperation from BRepAlgoAPI; 
    ---Purpose:  Empty constructor   
    -- <PF> - PaveFiller object that is carried out  
     
    Initialize (S1 :Shape from TopoDS;  
                S2 :Shape from TopoDS; 
                anOperation:Operation from BOPAlgo); 
    ---Purpose: Constructor with two arguments  
    -- <S1>, <S2>  -arguments     
    -- <anOperation> - the type of the operation
    -- Obsolete 
     
    Initialize (S1 :Shape from TopoDS; 
                S2 :Shape from TopoDS; 
                PF :PaveFiller from BOPAlgo;               
                anOperation:Operation from BOPAlgo); 
    ---Purpose: Constructor with two arguments  
    -- <S1>, <S2>  -arguments     
    -- <anOperation> - the type of the operation 
    -- <PF> - PaveFiller object that is carried out  
    -- Obsolete  
    
    Shape1(me)   
        returns Shape from TopoDS 
        is static; 
    ---Purpose: Returns the first argument involved in this Boolean operation. 
    -- Obsolete 
    ---C++: return const &
    

    Shape2(me)  
        returns Shape from TopoDS 
        is static;
    ---Purpose: Returns the second argument involved in this Boolean operation. 
    -- Obsolete 
    ---C++: return const &
      
    SetTools(me:out; 
           theLS: ListOfShape from BOPCol); 
    ---Purpose: Sets the tools    
     
    Tools(me) 
      returns ListOfShape from BOPCol; 
    ---C++: return const &   
    ---Purpose: Gets the tools    
     
    SetOperation (me:out; 
            anOp:  Operation from BOPAlgo);  
    ---Purpose:  Sets the type of Boolean operation 
     
    Operation  (me) 
        returns Operation from BOPAlgo;
    ---Purpose: Returns the type of Boolean Operation 
    ---C++: alias "Standard_EXPORT virtual ~BRepAlgoAPI_BooleanOperation();"  
    
    Build  (me:out) 
        is redefined ; 
    ---Purpose: Performs the algorithm 
    -- Filling interference Data Structure (if it is necessary)
    -- Building the result of the operation. 
     
    BuilderCanWork(me)  
        returns Boolean from Standard;  
    ---Purpose: Returns True if there was no errors occured 
    -- obsolete 
     
    FuseEdges(me)   
        returns Boolean from Standard;
    ---Purpose: Returns the flag of edge refining  
     
    RefineEdges(me:out);
    ---Purpose: Fuse C1 edges
     
    SectionEdges (me:  in  out)  
        returns ListOfShape from TopTools;    
    --- Purpose: Returns a list of section edges.
    -- The edges represent the result of intersection between arguments of
    -- Boolean Operation. They are computed during operation execution.
    ---C++:  return const &  
         
    Modified (me: in out;  
            aS : Shape from TopoDS) 
        returns ListOfShape from TopTools
        is redefined;
    ---Purpose: Returns the list  of shapes modified from the shape <S>. 
    ---C++: return const & 

    IsDeleted (me: in out;  
            aS : Shape from TopoDS)
        returns Boolean
        is redefined;
    ---Purpose: Returns true if the shape S has been deleted. The
    -- result shape of the operation does not contain the shape S.
        
    Generated (me: in out;  
            S : Shape from TopoDS)
        returns ListOfShape from TopTools
        is redefined;
    ---Purpose: Returns the list  of shapes generated from the shape <S>.
    ---         For use in BRepNaming.
    ---C++:  return const &
    
    HasModified (me) 
        returns Boolean from Standard
        is redefined;
    ---Purpose: Returns true if there is at least one modified shape.
    ---         For use in BRepNaming.

    HasGenerated (me)
        returns Boolean from Standard
        is redefined;
    ---Purpose: Returns true if there is at least one generated shape.
    ---         For use in BRepNaming.

    HasDeleted (me)
        returns Boolean from Standard
        is redefined;
    ---Purpose: Returns true if there is at least one deleted shape.
    ---         For use in BRepNaming.
 
    --  
    -- protected methods
    --     
    Clear(me:out) 
        is redefined protected;  
	 
    SetAttributes (me:out) 
        is virtual protected;   
	
    RefinedList (me:  in  out;  
            theL : ListOfShape from TopTools)  
        returns ListOfShape from TopTools
        is protected;
    ---Purpose: Returns the list  of shapes generated from the shape <S>.
    ---         For use in BRepNaming.
    ---C++:  return const & 
     
    
    
fields 
    myTools    : ListOfShape from BOPCol is protected; 
    myOperation: Operation from BOPAlgo   is protected;   
    -- 
    myBuilderCanWork : Boolean from Standard is protected;   
    --    for  edge  refiner
    myFuseEdges      : Boolean from Standard ; 
    myModifFaces     : DataMapOfShapeShape from TopTools;   
    myEdgeMap        : DataMapOfShapeShape from TopTools; 
    
end BooleanOperation;
