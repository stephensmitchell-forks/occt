-- Created on: 1994-07-12
-- Created by: Bruno DUMORTIER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakePipe from BRepOffsetAPI inherits MakeSweep from BRepPrimAPI

    	---Purpose: Describes functions to build pipes.
    	-- A pipe is built a basis shape (called the profile) along
    	-- a wire (called the spine) by sweeping.
    	-- The profile must not contain solids.
    	-- A MakePipe object provides a framework for:
    	-- - defining the construction of a pipe,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result.
    	-- Warning
    	-- The MakePipe class implements pipe constructions
    	-- with G1 continuous spines only.
uses
    Pipe        from BRepFill,
    Trihedron   from GeomFill,
    Wire        from TopoDS,
    Shape       from TopoDS,
    Edge        from TopoDS,
    ListOfShape from TopTools

is


    Create( Spine   : Wire  from TopoDS;
    	    Profile : Shape from TopoDS )
	---Purpose: Constructs a pipe by sweeping the shape Profile along
    	-- the wire Spine.The angle made by the spine with the profile is
    	-- maintained along the length of the pipe.
    	-- Warning
    	-- Spine must be G1 continuous; that is, on the connection
    	-- vertex of two edges of the wire, the tangent vectors on
    	-- the left and on the right must have the same direction,
    	-- though not necessarily the same magnitude.
        -- Exceptions
    	-- Standard_DomainError if the profile is a solid or a
    	-- composite solid.
    returns MakePipe from BRepOffsetAPI;

    Create( Spine   : Wire  from TopoDS;
    	    Profile : Shape from TopoDS;
	    aMode   : Trihedron from GeomFill;
	    ForceApproxC1 : Boolean from Standard = Standard_False)
	---Purpose: the same as previous but with setting of
	--          mode of sweep and the flag that indicates attempt
	--          to approximate a C1-continuous surface if a swept
	--          surface proved to be C0.
    returns MakePipe from BRepOffsetAPI;

    Pipe(me) returns Pipe from BRepFill
	---C++: return const &
	---Level: Advanced
    is static;


    Build(me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeShape).
	---Level: Public


    FirstShape (me : in out)
    ---Purpose: Returns the  TopoDS  Shape of the bottom of the prism.
    returns Shape from TopoDS;


    LastShape (me : in out)
    ---Purpose: Returns the TopoDS Shape of the top of the prism.
    returns Shape from TopoDS;

    Generated (me: in out; S: Shape from TopoDS)
    returns ListOfShape from TopTools
    is redefined;
    ---C++: return const &
    ---Level: Public

    Generated (me: in out; SSpine, SProfile : Shape from TopoDS)
        ---Level: Public
    returns Shape from TopoDS;


    ErrorOnSurface (me)
        ---Level: Public
    returns Real from Standard;


fields

    myPipe : Pipe from BRepFill;

end MakePipe;
