-- Created on: 2004-01-09
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class GeomTolerance from XCAFDoc inherits Attribute from TDF

	---Purpose: attribute to store dimension and tolerance

uses
    Label from TDF,
    RelocationTable from TDF,
    GeomToleranceObject from XCAFDimTolObjects

is

    Create returns GeomTolerance from XCAFDoc;

    Create(theObj : GeomTolerance from XCAFDoc) returns GeomTolerance from XCAFDoc;
    
    ---Category: class methods
    --           =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;

    Set (myclass; theLabel : Label from TDF)
    returns GeomTolerance from XCAFDoc;

    SetObject (me : mutable; theObject : GeomToleranceObject from XCAFDimTolObjects);

    GetObject (me) returns GeomToleranceObject from XCAFDimTolObjects;
                                                                                
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    


end GeomTolerance;
