-- Created by: Peter KURNEV
-- Copyright (c) 2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class BuilderAlgo from BRepAlgoAPI
        inherits Algo from BRepAlgoAPI 
    ---Purpose:  
    --  The clsss contains API level of General Fuse algorithm

uses
    Shape from TopoDS, 
    ListOfShape from TopTools,
    ListOfShape from BOPCol,
    --
    PPaveFiller from BOPAlgo, 
    PaveFiller from BOPAlgo,
    PBuilder from BOPAlgo
    
--raises

is
    Create  
        returns BuilderAlgo from BRepAlgoAPI; 
    ---Purpose:  Empty constructor 
    ---C++: alias "Standard_EXPORT virtual ~BRepAlgoAPI_BuilderAlgo();"

 
    Create(thePF  :PaveFiller from BOPAlgo)  
        returns BuilderAlgo from BRepAlgoAPI; 
    ---Purpose:  Empty constructor  
     
    SetFuzzyValue(me:out; 
        theFuzz : Real from Standard);
    ---Purpose: Sets the additional tolerance

    FuzzyValue(me)
        returns Real from Standard;
    ---Purpose: Returns the additional tolerance   
    
    SetArguments(me:out; 
        theLS: ListOfShape from BOPCol);  
    ---Purpose: Sets the arguments    
            
    Arguments(me) 
        returns ListOfShape from BOPCol; 
    ---C++: return const & 
    ---Purpose: Gets the arguments   
    
    Build  (me:out) 
        is redefined virtual; 
    ---Purpose:  Performs the algorithm 
    -- 
    --  H  I  S  T  O  R  Y           
    --
    Modified (me: in out;  
            aS : Shape from TopoDS) 
        returns ListOfShape from TopTools
        is redefined virtual;
    ---Purpose: Returns the list  of shapes modified from the shape <S>. 
    ---C++: return const & 

    IsDeleted (me: in out;  
            aS : Shape from TopoDS)
        returns Boolean
        is redefined virtual;
    ---Purpose: Returns true if the shape S has been deleted. The
    -- result shape of the operation does not contain the shape S.
        
    Generated (me: in out;  
            S : Shape from TopoDS)
        returns ListOfShape from TopTools
        is redefined virtual;
    ---Purpose: Returns the list  of shapes generated from the shape <S>.
    ---         For use in BRepNaming.
    ---C++:  return const &
    
    HasModified (me) 
        returns Boolean from Standard
        is virtual;
    ---Purpose: Returns true if there is at least one modified shape.
    ---         For use in BRepNaming.

    HasGenerated (me)
        returns Boolean from Standard
        is virtual;
    ---Purpose: Returns true if there is at least one generated shape.
    ---         For use in BRepNaming.

    HasDeleted (me)
        returns Boolean from Standard
        is virtual;
    ---Purpose: Returns true if there is at least one deleted shape.
    ---         For use in BRepNaming. 
    --
    --  protected methods
    --
    Clear(me:out) 
        is redefined protected; 

fields
    myEntryType  : Integer from Standard is protected;    
    myDSFiller   : PPaveFiller from BOPAlgo  is protected;
    myBuilder    : PBuilder    from BOPAlgo  is protected;
    myFuzzyValue : Real        from Standard is protected; 
    myArguments  : ListOfShape from BOPCol is protected;   
end BuilderAlgo;
