-- Created on: 1997-12-18
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Reader from PCDM inherits Transient from Standard


uses
    Document from CDM, 
    ExtendedString from TCollection,  
    Application from CDM, 
    ReaderStatus from PCDM,
    IStream from Standard,
    Data from Storage
		      
raises  DriverError from PCDM


is

    CreateDocument(me: mutable) returns Document from CDM
    is deferred;
    ---Purpose: this method is called by the framework before the read method.
    
    Read(me: mutable; aFileName: ExtendedString from TCollection; 
                      aNewDocument: Document from CDM;
		      anApplication: Application from CDM)
    raises DriverError from PCDM
    is deferred;
    ---Purpose: retrieves the content of the file into a new Document.  

    Read(me: mutable; theIStream:  in out IStream from Standard;
                      theStorageData: Data from Storage;
                      aNewDocument: Document from CDM;
		      anApplication: Application from CDM)
    raises DriverError from PCDM
    is deferred;
    ---Purpose: retrieves the content of the stream into a new Document.  
    
    GetStatus(me) returns ReaderStatus from PCDM; 
    ---C++: inline
fields 

    myReaderStatus : ReaderStatus from  PCDM is protected;
    
end Reader from PCDM;

