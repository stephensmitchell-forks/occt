-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

deferred  class ModelModifier from IGESSelect inherits Modifier from IFSelect
uses CString,
     InterfaceModel,
     Protocol from Interface,
     Protocol from IGESData,
     IGESModel from IGESData,
     CopyTool from Interface,
     ContextModif

is
    Initialize(mayChangeGraph : Boolean);
    ---Purpose : Calls inherited Initialize, transmits to it the information
    --           <mayChangeGraph>

    Perform (me; theContext  : in out ContextModif from IFSelect;
    	     theTarget   : mutable InterfaceModel from Interface;
    	     theProtocol : Protocol from Interface;
    	     theCopyTool       : in out CopyTool from Interface);
    ---Purpose : The inherited Perform does the required cast (and refuses to
    --           go further if cast has failed) then calls the instantiated
    --           Performing

    PerformProtocol (me; theContext : in out ContextModif  from IFSelect;
    	     theTarget : mutable IGESModel from IGESData;
    	     theProtocol  : Protocol from IGESData;
    	     theCopyTool     : in out CopyTool from Interface)  is virtual;
    ---Purpose : Specific Perform with Protocol. It is defined to let the
    --           Protocol unused and to call Performing without Protocol
    --           (most current case). It can be redefined if specific action
    --           requires Protocol.

    Performing (me; theContext : in out ContextModif from IFSelect;
    	     theTarget : mutable IGESModel from IGESData;
    	     theCopyTool     : in out CopyTool from Interface)  is deferred;
    ---Purpose : Specific Perform, without Protocol. If Performing with
    --           Protocol is redefined, Performing without Protocol must
    --           though be defined to do nothing (not called, but demanded
    --           by the linker)

end ModelModifier;