-- Created on: 1994-03-22
-- Created by: Frederic UNTEREINER
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package IGESToBRep

    ---Purpose : Provides tools in order to transfer IGES entities
    --         to CAS.CADE.

uses

    Interface,
    Transfer,
    MoniTool,
    Message,
    IGESData,
    IGESBasic,
    IGESGeom,
    IGESSolid,
    gp,
    Geom,
    Geom2d,
    TColGeom,
    TColGeom2d,
    TColStd,
    TopoDS,
    TopTools,
    ShapeExtend,
    ShapeAnalysis
    
is

    class CurveAndSurface;
    	class BasicSurface;
    	class BasicCurve;
    	class TopoSurface;
    	class TopoCurve;
    	class BRepEntity;

    class IGESBoundary;
    imported Reader;
    imported Actor;
    class AlgoContainer;
    class ToolContainer;
 
    Init;                                                                                                                
        ---Purpose: Creates and initializes default AlgoContainer.     
 
    SetAlgoContainer (aContainer: AlgoContainer from IGESToBRep);                                                          
        ---Purpose: Sets default AlgoContainer                                                                           
                                                                                                                         
    AlgoContainer returns AlgoContainer from IGESToBRep;                                                                   
        ---Purpose: Returns default AlgoContainer    
	
    IsCurveAndSurface(start : IGESEntity from IGESData)
    	returns Boolean;
        ---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferCurveAndSurface.
    	--          ex: All IGESEntity from IGESGeom


    IsBasicCurve  (start : IGESEntity from IGESData)
    	returns Boolean;
    	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferBasicCurve.
    	--          ex: CircularArc, ConicArc, Line, CopiousData,
    	--              BSplineCurve, SplineCurve... from IGESGeom :
    	--              104,110,112,126


    IsBasicSurface(start : IGESEntity from IGESData)
    	returns Boolean;
      	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferBasicSurface.
    	--          ex: BSplineSurface, SplineSurface... from IGESGeom :
    	--              114,128
     

    IsTopoCurve(start : IGESEntity from IGESData)
    	returns Boolean;
      	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferTopoCurve.         
    	--          ex: all Curves from IGESGeom :
    	--              all basic curves,102,130,142,144

     
    IsTopoSurface(start : IGESEntity from IGESData)
    	returns Boolean;
     	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferTopoSurface.
    	--          ex: All Surfaces from IGESGeom : 
    	--              all basic surfaces,108,118,120,122,141,143
     

    IsBRepEntity  (start : IGESEntity from IGESData)
    	returns Boolean;
    	---Purpose: Return True if the IGESEntity can be transfered by
    	--          TransferBRepEntity.
    	--          ex: VertexList, EdgeList, Loop, Face, Shell, 
    	--              Manifold Solid BRep Object from IGESSolid :
    	--              502, 504, 508, 510, 514, 186.

    WriteShape(shape  : Shape from TopoDS;
    	       number : Integer from Standard);
    	---Purpose: Creates  a file  Shape_'number' with the shape being
    	--          able to be restored by Draw.

    IGESCurveToSequenceOfIGESCurve (curve   : IGESEntity from IGESData;
    	    	    	    	    sequence: out HSequenceOfTransient from TColStd)
    returns Integer;
    
    TransferPCurve (fromedge: Edge from TopoDS;
    	    	    toedge  : Edge from TopoDS;
    	    	    face    : Face from TopoDS)
    returns Boolean;
    
end IGESToBRep;


