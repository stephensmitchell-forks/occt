-- Created on: 1993-10-14
-- Created by: Remi LEQUETTE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Fuse from BRepAlgoAPI inherits BooleanOperation from BRepAlgoAPI

        ---Purpose:  The class Fuse provides a
            -- Boolean fusion operation on a pair of arguments (Boolean Union).
            -- The class Fuse provides a framework for:
            --   -       Defining the construction of a fused shape;
            --   -       Implementing the building algorithm
            --   -       Consulting the result.

uses
    Shape from TopoDS, 
    PaveFiller from BOPAlgo

is
    Create (S1, S2  : Shape from TopoDS; 
            theFuzz : Real from Standard = 0.0)  
            returns Fuse from BRepAlgoAPI;  
        ---Purpose: Constructs a fuse of shapes aS1 and aS2.
         
    Create (S1,S2 : Shape from TopoDS; 
            aDSF  : PaveFiller from BOPAlgo)  
            returns Fuse from BRepAlgoAPI; 
        ---Purpose: Constructs a new shape that is a fuse of shapes aS1 and aS2 using aDSFiller. 
    
end Fuse;
