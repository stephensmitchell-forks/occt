-- Created on: 1997-12-09
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

private class ReadWriter_1 from PCDM inherits ReadWriter from PCDM

uses
    ExtendedString from TCollection,  
    AsciiString from TCollection, 
    Data from Storage, 
    IODevice from Storage,
    Document from CDM, 
    MessageDriver from CDM, 
    SequenceOfExtendedString from TColStd, 
    SequenceOfReference from PCDM

is

    Create returns ReadWriter_1 from PCDM;
   
    Version(me) returns AsciiString from TCollection;
    ---Purpose: returns PCDM_ReadWriter_1.
   
    WriteReferenceCounter(me; aData: Data from Storage; aDocument: Document from CDM);

    WriteReferences(me; aData: Data from Storage; aDocument: Document from CDM; theReferencer: IODevice from Storage);

    WriteExtensions(me; aData: Data from Storage; aDocument: Document from CDM);

    WriteVersion(me; aData: Data from Storage; aDocument: Document from CDM);
    
    ReadReferenceCounter(me; aDevice: IODevice from Storage; theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard;

    ReadReferences(me; aDevice: IODevice from Storage; theReferences: in out  SequenceOfReference from PCDM; theMsgDriver: MessageDriver from CDM);

    
    ReadExtensions(me; aDevice: IODevice from Storage; theExtensions: in out  SequenceOfExtendedString from TColStd; theMsgDriver: MessageDriver from CDM);

    ReadUserInfo(myclass; aDevice: IODevice from Storage; Start, End: AsciiString from TCollection; theUserInfo:in  out SequenceOfExtendedString from TColStd;theMsgDriver: MessageDriver from CDM)
    is private;

    ReadDocumentVersion(me; aDevice: IODevice from Storage; theMsgDriver: MessageDriver from CDM)
    returns Integer from Standard;

end ReadWriter_1 from PCDM;
