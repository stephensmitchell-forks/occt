---Copyright: Open CASCADE 2014
-- Created on: 2012-06-09
-- Created by: jgv@ROLEX
-- Copyright (c) 2012-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class UnifySameDomain from ShapeUpgrade inherits TShared from MMgt

	---Purpose: Unifies same domain faces and edges of specified shape

uses
    Shape from TopoDS,
    ListOfShape from TopTools,
    DataMapOfShapeShape from TopTools,
    ReShape from ShapeBuild

is
    Create returns UnifySameDomain from ShapeUpgrade;
    ---Purpose: empty constructor

    Create(aShape: Shape from TopoDS;
    	   UnifyEdges: Boolean from Standard = Standard_True;
	   UnifyFaces: Boolean from Standard = Standard_True;
    	   ConcatBSplines: Boolean from Standard = Standard_False)
    returns UnifySameDomain from ShapeUpgrade;
    
    Initialize(me: mutable; aShape: Shape from TopoDS;
    	       UnifyEdges: Boolean from Standard = Standard_True;
	       UnifyFaces: Boolean from Standard = Standard_True;
    	       ConcatBSplines: Boolean from Standard = Standard_False);
    
    Build( me : mutable );
    	---Purpose: Builds the resulting shape
    
    Shape(me) returns Shape from TopoDS;
    	---C++: return const &
    	---Purpose: Gives the resulting shape
    
    Generated (me; aShape : Shape from TopoDS)
    returns Shape from TopoDS;
    
    UnifyFaces(me: mutable);
    ---Purpose: this method makes if possible a common face from each
    --          group of faces lying on coincident surfaces

    UnifyEdges(me: mutable);
    ---Purpose: this method makes if possible a common edge from each
    --          group of edges connecting common couple of faces

    UnifyFacesAndEdges(me: mutable);
    ---Purpose: this method unifies same domain faces and edges

fields
    
    myInitShape : Shape from TopoDS;
    myUnifyFaces : Boolean from Standard;
    myUnifyEdges : Boolean from Standard;
    myConcatBSplines : Boolean from Standard;
    
    myShape : Shape from TopoDS;
    
    myContext   : ReShape from ShapeBuild;
    myOldShapes : DataMapOfShapeShape from TopTools;
    
end UnifySameDomain;
