-- Created on: 1994-12-22
-- Created by: Christian CAILLET
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package StepSelect

    ---Purpose : This package defines the library of the tools used for every
    --           kind of STEP Files, i.e. whatever the considered Protocol.

uses MMgt, TCollection, TColStd, Message,
     Interface, IFGraph, IFSelect, StepData

is

    class StepType;

    imported FileModifier;

    imported FloatFormat;

    class WorkLibrary;

    class Activator;

end StepSelect;
