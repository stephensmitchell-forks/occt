-- Created on: 2001-07-25
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2001-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XmlLDrivers

uses
    Standard,
    Storage,
    TDF,
    TDocStd,
    TCollection,
    TColStd,
    CDM,
    PCDM,
    XmlObjMgt,
    XmlMDF

is
    class DocumentStorageDriver;
    class DocumentRetrievalDriver;

    private class NamespaceDef;
    
    private class SequenceOfNamespaceDef
        instantiates Sequence from TCollection (NamespaceDef from XmlLDrivers);

    Factory (theGUID : GUID from Standard) returns Transient from Standard;

    CreationDate returns AsciiString from TCollection;

    AttributeDrivers (theMsgDriver: MessageDriver from CDM)
        returns ADriverTable from XmlMDF; 
	
    StorageVersion returns AsciiString from TCollection; 
    
end XmlLDrivers;
