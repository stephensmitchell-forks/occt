-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class Algo from BOPAlgo 
	---Purpose: provides the root interface for algorithms

uses  
    BaseAllocator from BOPCol

--raises

is
    Initialize 
    	returns Algo from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_Algo();"  
     
    Initialize (theAllocator: BaseAllocator from BOPCol) 
    	returns Algo from BOPAlgo;  
     
    Perform(me:out) 
	is deferred;      
         
    ErrorStatus (me) 
    	returns Integer from Standard; 
  
    WarningStatus (me) 
    	returns Integer from Standard;
  
    CheckData(me:out) 
	is virtual protected;  
    	
    CheckResult(me:out) 
	is virtual protected; 

    Allocator(me) 
    	returns BaseAllocator from BOPCol; 
    ---C++: return const &	
 
    SetRunParallel(me:out; 
    	    theFlag:Boolean from Standard); 
    ---Purpose: Set the flag of parallel processing 
    -- if <theFlag> is true  the parallel processing is switched on   
    -- if <theFlag> is false the parallel processing is switched off   
    --      
    RunParallel(me) 
    	returns Boolean from Standard; 
    ---Purpose: Returns the flag of parallel processing  

fields 
    myAllocator     : BaseAllocator from BOPCol is protected;
    myErrorStatus   : Integer from Standard is protected;	 
    myWarningStatus : Integer from Standard is protected;	 
    myRunParallel : Boolean from Standard is protected; 
end Algo;
