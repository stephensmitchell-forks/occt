-- Created on: 1999-09-08
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ValidationProps from STEPConstruct inherits Tool from STEPConstruct

    ---Purpose: This class provides tools for access (write and read)
    --          the validation properties on shapes in the STEP file.
    --          These are surface area, solid volume and centroid.

uses
    WorkSession_Handle        from XSControl,
    InterfaceModel     from Interface,
    HGraph             from Interface,
    FinderProcess_Handle      from Transfer,
    TransientProcess_Handle   from Transfer,
    RepresentationItem from StepRepr,
    Pnt                from gp,
    Shape              from TopoDS,
    MapOfShape         from TopTools,
    SequenceOfTransient from TColStd,
    Unit                from StepBasic,
    CharacterizedDefinition from StepRepr,
    RepresentationContext from StepRepr,
    --ShapeDefinitionRepresentation from StepShape,
    --ContextDependentShapeRepresentation from StepShape,
    ProductDefinition     from StepBasic,
    NextAssemblyUsageOccurrence from StepRepr,
    PropertyDefinition    from StepRepr,
    RepresentationContext from StepRepr

is

    Create returns ValidationProps;
    	---Purpose: Creates an empty tool

    Create (WS: WorkSession_Handle from XSControl) returns ValidationProps;
    	---Purpose: Creates a tool and loads it with worksession
	
    Init (me: in out; WS: WorkSession_Handle from XSControl) returns Boolean;
    	---Purpose: Load worksession; returns True if succeeded
	
    AddProp (me: in out; Shape: Shape from TopoDS; 
                         Prop: RepresentationItem from StepRepr;
    	    	    	 Descr: CString;
    	    	    	 instance: Boolean = Standard_False)
    returns Boolean;
	---Purpose: General method for adding (writing) a validation property 
	--          for shape which should be already mapped on writing itself.
	--          It uses FindTarget() to find target STEP entity
        --          resulting from given shape, and associated context
	--          Returns True if success, False in case of fail
	
    AddProp (me: in out; target: CharacterizedDefinition from StepRepr;
    	    	    	 Context: RepresentationContext from StepRepr;
    	    	    	 Prop: RepresentationItem from StepRepr;
    	    	    	 Descr: CString)
    returns Boolean;
	---Purpose: General method for adding (writing) a validation property 
	--          for shape which should be already mapped on writing itself.
	--          It takes target and Context entities which correspond to shape
	--          Returns True if success, False in case of fail
	
							 
    AddArea (me: in out; Shape: Shape from TopoDS; Area: Real)
    returns Boolean;
        ---Purpose: Adds surface area property for given shape (already mapped).
	--          Returns True if success, False in case of fail

    AddVolume (me: in out; Shape: Shape from TopoDS; Vol: Real)
    returns Boolean;
        ---Purpose: Adds volume property for given shape (already mapped).
	--          Returns True if success, False in case of fail

    AddCentroid (me: in out; Shape: Shape from TopoDS; Pnt: Pnt from gp;
    	    	    	     instance: Boolean = Standard_False)
    returns Boolean;
        ---Purpose: Adds centroid property for given shape (already mapped).
	--          Returns True if success, False in case of fail
	--          If instance is True, then centroid is assigned to
	--          an instance of component in assembly

    FindTarget (me: in out; S: Shape from TopoDS;
    	    	    	    target: out CharacterizedDefinition from StepRepr;
    	    	    	    Context: out RepresentationContext from StepRepr;
    	    	    	    instance: Boolean = Standard_False)
    returns Boolean;
	---Purpose: Finds target STEP entity to which validation props should
	--          be assigned, and corresponding context, starting from shape
	--          Returns True if success, False in case of fail
	
    LoadProps (me; seq: out SequenceOfTransient from TColStd) returns Boolean;
    	---Purpose: Searches for entities of the type PropertyDefinitionRepresentation
	--          in the model and fills the sequence by them
	
    GetPropNAUO (me; PD: PropertyDefinition from StepRepr)
    returns     NextAssemblyUsageOccurrence from StepRepr;
    	---Purpose: Returns CDSR associated with given PpD or NULL if not found
	--          (when, try GetPropSDR)
	
    GetPropPD (me; PD: PropertyDefinition from StepRepr)
    returns ProductDefinition from StepBasic;
    	---Purpose: Returns SDR associated with given PpD or NULL if not found
	--          (when, try GetPropCDSR)
	
    GetPropShape (me; ProdDef: ProductDefinition from StepBasic)
    returns Shape from TopoDS;
    	---Purpose: Returns Shape associated with given SDR or Null Shape 
	--          if not found
    
    GetPropShape (me; PD: PropertyDefinition from StepRepr)
    returns Shape from TopoDS;
    	---Purpose: Returns Shape associated with given PpD or Null Shape 
	--          if not found
	
    GetPropReal (me; item: RepresentationItem from StepRepr; 
    	    	     Val: out Real; isArea: out Boolean)
    returns Boolean;
    	---Purpose: Returns value of Real-Valued property (Area or Volume)
	--          If Property is neither Area nor Volume, returns False
	--          Else returns True and isArea indicates whether property
	--          is area or volume
	
    GetPropPnt (me; item: RepresentationItem from StepRepr; 
    	    	    Context: RepresentationContext from StepRepr;
    	    	    Pnt: out Pnt from gp)
    returns Boolean;
    	---Purpose: Returns value of Centriod property (or False if it is not)
	
    SetAssemblyShape (me: in out; shape: Shape from TopoDS);
    	---Purpose: Sets current assembly shape SDR (for FindCDSR calls)
	
fields

    areaUnit, volUnit: Unit from StepBasic; -- units for sharing on writing
    myAssemblyPD: ProductDefinition from StepBasic;

end ValidationProps;
