-- Created on: 2004-01-15
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Datum from XCAFDoc inherits Attribute from TDF

	---Purpose: attribute to store datum

uses
    Label from TDF,
    RelocationTable from TDF,
    HAsciiString from TCollection,
    DatumObject from XCAFDimTolObjects

is
 
    Create returns Datum from XCAFDoc;
    
    ---Category: class methods
    --           =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;
    
    Set (myclass; label : Label from TDF;
    	    	  aName : HAsciiString from TCollection;
    	    	  aDescription : HAsciiString from TCollection;
    	    	  anIdentification : HAsciiString from TCollection)
    returns Datum from XCAFDoc;

    Set (myclass; label : Label from TDF)
    returns Datum from XCAFDoc;


    Set (me : mutable; aName : HAsciiString from TCollection;
    	    	       aDescription : HAsciiString from TCollection;
    	    	       anIdentification : HAsciiString from TCollection);
	     
    GetName (me) returns HAsciiString from TCollection;
                                                                   
    GetDescription (me) returns HAsciiString from TCollection;

    GetIdentification (me) returns HAsciiString from TCollection;

    GetObject (me) returns DatumObject from XCAFDimTolObjects;

    SetObject (me : mutable; theObject : DatumObject from XCAFDimTolObjects);

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

fields
    myName : HAsciiString from TCollection;
    myDescription : HAsciiString from TCollection;
    myIdentification : HAsciiString from TCollection;

end Datum;
