-- Created on: 1993-01-13
-- Created by: CKY / Contract Toubro-Larsen ( Deepak PRABHU )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class AssociativityDef from IGESDefs  inherits IGESEntity

        ---Purpose: defines IGES Associativity Definition Entity, Type <302>
        --          Form <5001 - 9999> in package IGESDefs.
        --          This class permits the preprocessor to define an
        --          associativity schema. i.e., by using it preprocessor
        --          defines the type of relationship.

uses

        HArray1OfInteger                 from TColStd,
        HArray1OfHArray1OfInteger_Handle from IGESBasic

raises DimensionMismatch, OutOfRange

is

        Create returns mutable AssociativityDef;

        -- Specific methods for the entity

        Init (me           : mutable;
              requirements : HArray1OfInteger;
              orders       : HArray1OfInteger;
              numItems     : HArray1OfInteger;
              items        : HArray1OfHArray1OfInteger_Handle)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           AssociativityDef
        --       - requirements : Back Pointers requirements
        --       - orders       : Class Orders
        --       - numItems     : Number of Items per Class
        --       - items        : Items in each class
        -- raises exception if lengths of the arrays are not the same.

    	SetFormNumber (me : mutable; form : Integer);
	-- Sets Form Number to a given value (free over 5000)


        NbClassDefs(me) returns Integer;
        ---Purpose : returns the Number of class definitions

        IsBackPointerReq(me ; ClassNum : Integer) returns Boolean
        raises OutOfRange;
        ---Purpose : returns 1 if the theBackPointerReqs(ClassNum) = 1
        -- returns 0 if the theBackPointerReqs(ClassNum) = 2
        -- raises exception if ClassNum <= 0 or ClassNum > NbClassDefs()

        BackPointerReq(me ; ClassNum : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns 1 or 2
        -- raises exception if ClassNum <= 0 or ClassNum > NbClassDefs()

        IsOrdered(me ; ClassNum : Integer) returns Boolean
        raises OutOfRange;
        ---Purpose : returns 1 if theClassOrders(ClassNum) = 1 (ordered class)
        -- returns 0 if theClassOrders(ClassNum) = 2 (unordered class)
        -- raises exception if ClassNum <= 0 or ClassNum > NbClassDefs()

        ClassOrder(me ; ClassNum : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns 1 or 2
        -- raises exception if ClassNum <= 0 or ClassNum > NbClassDefs()

        NbItemsPerClass(me ; ClassNum : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns no. of items per class entry
        -- raises exception if ClassNum <= 0 or ClassNum > NbClassDefs()

        Item(me ; ClassNum : Integer; ItemNum : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns ItemNum'th Item of ClassNum'th Class
        -- raises exception if
        --      ClassNum <= 0 or ClassNum > NbClassDefs()
        --      ItemNum <= 0 or ItemNum > NbItemsPerClass(ClassNum)

fields

--
--  Class    : IGESDefs_AssociativityDef
--
--  Purpose  : Declaration of variables specific to AssociativityDef
--
--  Reminder : An AssociativityDef Entity permits the preprocessor
--             to define an associativity schema. The definition
--             includes associativity form, the no. of classes,
--             the number and type of items in each class, and
--             whether back pointers are required.

        theBackPointerReqs : HArray1OfInteger;
        theClassOrders     : HArray1OfInteger;
        theNbItemsPerClass : HArray1OfInteger;
        theItems           : HArray1OfHArray1OfInteger_Handle;

end AssociativityDef;
