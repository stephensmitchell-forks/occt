-- Created on: 1994-07-06
-- Created by: Laurent PAINNOT
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class ExtCC from Extrema

    ---Purpose: It calculates all the distance between two curves.
    --          These distances can be maximum or minimum.

uses POnCurv           from Extrema,
     SequenceOfPOnCurv from Extrema,
     ExtElC            from Extrema,
     Pnt               from gp,
     HArray1OfPnt      from TColgp,
     SequenceOfReal    from TColStd,
     ListOfTransient   from TColStd,
     Curve             from Adaptor3d,
     CurveTool         from Extrema,
     ECC               from Extrema


raises  InfiniteSolutions from StdFail,
        NotDone           from StdFail,
        OutOfRange        from Standard


is

    Create (TolC1: Real = 1.0e-10; TolC2: Real = 1.0e-10) returns ExtCC;
    

    Create (C1: Curve from Adaptor3d;  C2: Curve from Adaptor3d;
            TolC1: Real = 1.0e-10; TolC2: Real = 1.0e-10) returns ExtCC;
      	---Purpose: It calculates all the distances.


    Create (C1: Curve from Adaptor3d;
    	    C2: Curve from Adaptor3d;
	    U1: Real  from Standard;
	    U2: Real  from Standard;
	    V1: Real  from Standard;
	    V2: Real  from Standard;
            TolC1: Real = 1.0e-10;
            TolC2: Real = 1.0e-10) returns ExtCC;
      	---Purpose: It calculates all the distances.


    SetCurve (me: in out; theRank: Integer; C: Curve from Adaptor3d);
        ---Purpose:

    SetCurve (me: in out; theRank: Integer; C: Curve from Adaptor3d; Uinf, Usup: Real);
        ---Purpose:

    SetRange (me: in out; theRank: Integer; Uinf, Usup: Real);
        ---Purpose:

    SetTolerance (me: in out; theRank: Integer; Tol: Real);
        ---Purpose:

    Perform(me: in out);
    

    IsDone (me) returns Boolean
    	---Purpose: Returns True if the distances are found.
    	is static;

    NbExt (me) returns Integer
    	---Purpose: Returns the number of extremum distances.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail
		-- if IsParallel(me)= True.
    	is static;


    IsParallel (me) returns Boolean
    	---Purpose: Returns True if the two curves are parallel.
    	raises  NotDone from StdFail
	    	-- if IsDone(me)=False.
    	is static;


    SquareDistance (me; N: Integer =1) returns Real
    	---Purpose: Returns the value of the Nth extremum square distance.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail,
		-- if IsParallel(me)= True and N > 1.
    	    	OutOfRange
		-- if N < 1 or N > NbExt(me)
    	is static;

    Points (me; N: Integer; P1,P2: out POnCurv)
    	---Purpose: Returns the points of the Nth extremum distance.
    	--          P1 is on the first curve, P2 on the second one.
    	raises  NotDone from StdFail,
	    	-- if IsDone(me)=False.
    	    	InfiniteSolutions from StdFail,
		-- if IsParallel(me)= True.
    	    	OutOfRange
		-- if N < 1 or N > NbExt(me)
    	is static;

    TrimmedSquareDistances(me; dist11, distP12, distP21, distP22: out Real;
                     P11, P12, P21, P22: out Pnt)
    	---Purpose: if the curve is a trimmed curve,
    	--          dist11 is a square distance between the point on C1
    	--          of parameter FirstParameter and the point of 
    	--          parameter FirstParameter on C2.

    is static;
    
    Results(me: in out; AlgExt: ExtElC from Extrema;
    	    Ut11, Ut12, Ut21, Ut22: Real)

    is static protected;    	

    Results(me: in out;AlgExt: ECC from Extrema;
    	    Ut11, Ut12, Ut21, Ut22: Real)

    is static protected;
    
    GetSingleSolutionFlag (me) returns Boolean
    ---Purpose: Returns single solution flag value.
    is static;
    
    SetSingleSolutionFlag (me: in out;
                           theFlag: Boolean)
    ---Purpose: Sets single solution flag value.
    is static;


    

fields
    myECC:    ECC from Extrema;
    myDone:   Boolean;
    myIsPar:  Boolean;
    myIsFindSingleSolution: Boolean;
    mypoints: SequenceOfPOnCurv from Extrema;
    mySqDist: SequenceOfReal    from TColStd;
    mynbext:  Integer;
    inverse:  Boolean;
    myC:     Address from Standard [2];
    myInf: Real [2];
    mySup: Real [2];
    myTol:  Real [2];
    P1f:      Pnt;
    P1l:      Pnt;
    P2f:      Pnt;
    P2l:      Pnt;
    mydist11: Real;
    mydist12: Real;
    mydist21: Real;
    mydist22: Real;
    


end ExtCC;
