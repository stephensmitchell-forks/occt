-- Created on: 1994-11-30
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MakeStepVertex from TopoDSToStep 
    inherits Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Vertex from TopoDS and TopologicalRepresentationItem from
    --          StepShape. 
  
uses Vertex                        from TopoDS,
     TopologicalRepresentationItem from StepShape,
     Tool                          from TopoDSToStep,
     MakeVertexError               from TopoDSToStep,
     FinderProcess_Handle                 from Transfer
          
raises NotDone from StdFail
     
is 

    Create returns MakeStepVertex;
    
    Create (V : Vertex from TopoDS;
    	    T : in out Tool from TopoDSToStep;
	   FP : FinderProcess_Handle from Transfer)
         returns MakeStepVertex;
    
    Init(me : in out;
     	 V  : Vertex from TopoDS;
     	 T  : in out Tool from TopoDSToStep;
         FP : FinderProcess_Handle from Transfer);

	    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const&
        
    Error(me) returns MakeVertexError from TopoDSToStep;

fields

    myResult : TopologicalRepresentationItem from StepShape;

    myError  : MakeVertexError from TopoDSToStep;
    
end MakeStepVertex;


