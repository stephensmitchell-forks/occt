-- Created on: 1995-01-25
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Presentation from PrsMgr
inherits TShared from MMgt

uses 

  PresentationManager from PrsMgr,
  NameOfColor from Quantity,
  Color       from Quantity,
  Transformation from Geom,
  Length from Quantity,
  ShadingAspect from Prs3d,
  TypeOfHighlightMethod from Aspect,
  TypeOfPresentation3d from PrsMgr,
  DataStructureManager from Graphic3d,
  Structure from Graphic3d,
  PresentableObjectPointer from PrsMgr,PresentableObject from PrsMgr,
  Prs from PrsMgr,
  Projector from Prs3d,
  Presentation from Prs3d

is

  Create (thePresentationManager : PresentationManager from PrsMgr;
          thePresentableObject   : PresentableObject   from PrsMgr)
  returns Presentation from PrsMgr
  is private;

  Destroy (me : mutable) is virtual;
  ---Level: Public
  ---Purpose: Destructor
  ---C++:     alias ~

  Display (me : mutable)
  is virtual private;

  Display (me : mutable;
           theIsHighlight : Boolean from Standard)
  is static private;
  ---Purpose: Displays myStructure.

  Erase (me : mutable)
  is virtual private;

  SetVisible (me       : mutable;
              theValue : Boolean from Standard)
  is virtual private;

  Highlight (me : mutable;
             theMethod : TypeOfHighlightMethod from Aspect;
             theColor  : Color                 from Quantity) is virtual private;

  Unhighlight (me) is virtual private;

  IsHighlighted (me) returns Boolean from Standard
  is virtual private;

  IsDisplayed (me) returns Boolean from Standard
  is virtual private;

  DisplayPriority(me) returns Integer from Standard
  is virtual private;

  SetDisplayPriority(me:mutable;aNewPrior:Integer from Standard)
  is virtual private;

  SetZLayer (me         : mutable;
             theLayerId : Integer from Standard)
  is virtual private;
  ---Purpose: Set Z layer ID for the presentation

  GetZLayer (me) returns Integer from Standard
  is virtual private;
  ---Purpose: Get Z layer ID for the presentation

  Clear (me : mutable)
  is virtual private;
  ---Purpose: removes the whole content of the presentation.
  --          Does not remove the other connected presentations.

---Category: references to other presentation.

  Connect (me;
           theOther : Presentation from PrsMgr)
  is static private;

---Category: Transformation methods.

  Transform (me;
             theTrsf : Transformation from Geom)
  is static private;

  Place (me;
         theX, theY, theZ : Length from Quantity)
  is static private;

  Multiply (me;
            theTrsf : Transformation from Geom)
  is static private;

  Move (me;
        theX, theY, theZ : Length from Quantity)
  is static private;

---Category: Global Aspect methods

  SetShadingAspect (me;
                    theShadingAspect : ShadingAspect from Prs3d)
  is static private;

  Presentation (me) returns Presentation from Prs3d
  is static;
  ---C++: inline
  ---C++: return const&

---Category: Computed Structures

  Compute (me           : mutable;
           theStructure : Structure from Graphic3d)
  is static private;

  Compute (me           : mutable;
           theProjector : DataStructureManager from Graphic3d)
  returns Structure from Graphic3d
  is static private;

  Compute (me           : mutable;
           theProjector : DataStructureManager from Graphic3d;
           theTrsf      : Transformation from Geom)
  returns Structure from Graphic3d
  is static private;

  Compute (me             : mutable;
           theProjector   : DataStructureManager from Graphic3d;
           theGivenStruct : Structure from Graphic3d)
  is static private;

  Compute (me             : mutable;
           theProjector   : DataStructureManager from Graphic3d;
           theTrsf        : Transformation from Geom;
           theGivenStruct : Structure from Graphic3d)
  is static private;

---Category: Inquire Methods

  PresentationManager (me) returns PresentationManager
  ---Purpose: returns the PresentationManager in which the presentation has been created.
  is static;
  ---C++: inline
  ---C++: return const&

  Projector (myclass;
             theProjector : DataStructureManager from Graphic3d)
  returns Projector from Prs3d
  is private;

---Category: Internal Methods

  SetUpdateStatus (me      : mutable;
                   theStat : Boolean from Standard);
  ---C++: inline

  MustBeUpdated (me) returns Boolean from Standard;
  ---C++: inline

fields

  myPresentationManager : PresentationManager from PrsMgr;
  myStructure           : Prs from PrsMgr;
  myPresentableObject   : PresentableObjectPointer from PrsMgr;
  myMustBeUpdated       : Boolean from Standard;
  myBeforeHighlightState: Integer from Standard;

friends

  class PresentationManager from PrsMgr,
  class PresentableObject   from PrsMgr,
  class Prs                 from PrsMgr

end Presentation from PrsMgr;
