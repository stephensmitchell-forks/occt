-- Created on: 1992-04-03
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PWalking from IntWalk
    
    ---Purpose: This class implements an algorithm to determine the
    --          intersection between 2 parametrized surfaces, marching from
    --          a starting point. The intersection line
    --          starts and ends on the natural surface's  boundaries .


uses XY                  from gp,
     StatusDeflection    from IntWalk,
     ConstIsoparametric  from IntImp,
     Array1OfReal        from TColStd,
     PntOn2S             from IntSurf,
     LineOn2S            from IntSurf,
     Dir                 from gp,
     Dir2d               from gp,
     Pnt                 from gp,
	 TheInt2S            from IntWalk,
     HSurface            from Adaptor3d,
     HSurfaceTool        from Adaptor3d
     
     
raises OutOfRange from Standard,
       NotDone    from StdFail
       

is


    Create ( Caro1 , 
             Caro2       : HSurface from Adaptor3d ; 
             TolTangency,
             Epsilon,
             Deflection,
             Increment   : Real from Standard)
	    
	---Purpose: Constructor used to set the data to compute intersection
	--          lines between Caro1 and Caro2.
    	--          Deflection is the maximum deflection admitted between two 
    	--          consecutive points on the resulting polyline.
    	--          TolTangency is the tolerance to find a tangent point.
    	--          Func is the criterion which has to be evaluated at each
    	--          solution point (each point of the line).
    	--          It is necessary to call the Perform method to compute 
    	--          the intersection lines.
    	--          The line found starts at a point on or in 2 natural domains
    	--          of surfaces. It can be closed in the 
    	--          standard case if it is open it stops and begins at the 
    	--          border of one of the domains. If an open line
    	--          stops at the middle of a domain, one stops at the tangent point.
    	--          Epsilon is SquareTolerance of points confusion.      

    	returns PWalking;
	

    Create ( Caro1 , 
             Caro2       : HSurface from Adaptor3d ; 
             TolTangency,
             Epsilon,
             Deflection,
             Increment   : Real from Standard;
             U1,V1,U2,V2 :Real from Standard)
	    
	---Purpose: Returns the intersection line containing the exact
	--          point Poin. This line is a polygonal line.
    	--          Deflection is the maximum deflection admitted between two 
    	--          consecutive points on the resulting polyline.
    	--          TolTangency is the tolerance to find a tangent point.
    	--          Func is the criterion which has to be evaluated at each
    	--          solution point (each point of the line).
    	--          The line found starts at a point on or in 2 natural domains
    	--          of surfaces. It can be closed in the 
    	--          standard case if it is open it stops and begins at the 
    	--          border of one of the domains. If an open line
    	--          stops at the middle of a domain, one stops at the tangent point.
    	--          Epsilon is SquareTolerance of points confusion.    

    	returns PWalking;

	
    Perform(me :in out;ParDep : Array1OfReal  from TColStd)
		       
    	---Purpose: calculate the line of intersection

    	is static;

    Perform(me :in out;ParDep : Array1OfReal  from TColStd;
    	    	u1min,v1min,u2min,v2min,u1max,v1max,u2max,v2max: Real from Standard)
		       
    	---Purpose: calculate the line of intersection. The regulation
    	--          of steps is done using min and max values on u and
    	--          v.  (if this data is not presented as in the
    	--          previous method, the initial steps are calculated
    	--          starting from min and max uv of faces).

    	is static;


    PerformFirstPoint(me :in out;
                      ParDep    : Array1OfReal  from TColStd;
                      FirstPoint: in out PntOn2S from IntSurf)
    
    	---Purpose: calculate the first point of a line of intersection
    	--          

    	returns Boolean from Standard

    	is static;


    IsDone(me)
    
    	---Purpose: Returns true if the calculus was successful.

    	returns Boolean from Standard
	---C++: inline

	is static;


    NbPoints(me)
    
    	---Purpose: Returns the number of points of the resulting polyline.
    	--          An exception is raised if IsDone returns False.

	returns Integer from Standard
	---C++: inline

	raises NotDone from StdFail

	is static;


    Value(me ; Index : Integer from Standard)
    
    	---Purpose: Returns the point of range Index on the polyline. 
    	--          An exception is raised if IsDone returns False.
    	--          An exception is raised if Index<=0 or Index>NbPoints.

    	returns  PntOn2S from IntSurf
	---C++: inline
	---C++: return const&

    	raises NotDone    from StdFail,
               OutOfRange from Standard
	
	is static;


    Line(me)
    
    	returns LineOn2S from IntSurf
	---C++: inline
	---C++: return const&
	
	raises NotDone from StdFail
	is static;


    TangentAtFirst(me)
    
    	---Purpose: Returns True if the surface are tangent at the first point
    	--          of the line.
    	--          An exception is raised if IsDone returns False.

    	returns Boolean from Standard
	---C++: inline

	raises NotDone from StdFail

	is static;


    TangentAtLast(me)
    
    	---Purpose: Returns true if the surface are tangent at the last point
    	--          of the line.
    	--          An exception is raised if IsDone returns False.

    	returns Boolean from Standard
	---C++: inline
	
	raises NotDone from StdFail
	is static;


    IsClosed(me)
    
    	---Purpose: Returns True if the line is closed.
    	--          An exception is raised if IsDone returns False.

	returns Boolean from Standard
	---C++: inline
	
	raises NotDone from StdFail
	is static;
      
      
    MaxStep(me ; Index : Integer from Standard)
    
    	---Purpose: Returns the point of range Index on the polyline. 
    	--          An exception is raised if IsDone returns False.
    	--          An exception is raised if Index<=0 or Index>NbPoints.

    	returns  Real from Standard
	---C++: inline

    	raises OutOfRange from Standard
	
	is static;
    	

    TangentAtLine(me; Index: out Integer from Standard)
    
    	returns Dir from gp
	---C++: return const&
	---C++: inline

	raises NotDone from StdFail
	is static;


--private

    TestDeflection(me : in out)

    	returns StatusDeflection from IntWalk
	is static;
	

    TestArret(me : in out; DejaReparti : Boolean from Standard;
                           Param : in out Array1OfReal from TColStd;
                           ChoixIso : out ConstIsoparametric from IntImp)


    	returns Boolean from Standard
	is static;
	

    RepartirOuDiviser(me : in out; DejaReparti : in out Boolean from Standard;
                      ChoixIso : out  ConstIsoparametric from IntImp;
		      Arrive : in out Boolean from Standard )
		      
	is static;

    AddAPoint ( me    : in out  ; 
    line  : in  out  LineOn2S  from  IntSurf  ;     
    POn2S :          PntOn2S   from  IntSurf  ) ;
    ---C++: inline
    
  ComputePasInit(me          : in out;
                 theDeltaU1, theDeltaV1, theDeltaU2, theDeltaV2: Real from Standard)

  is protected;

    
    ExtendLineInCommonZone(me: in out; theChoixIso: ConstIsoparametric  from IntImp;
theDirectionFlag: Boolean from Standard)
    returns Boolean from Standard
    is private;
  
  DistanceMinimizeByGradient( me    : in out;
                              theASurf1 , theASurf2  : HSurface from Adaptor3d ;
                              theU1, theV1, theU2, theV2: out Real from Standard;
                              theStep0U1V1: Real from Standard = 1.0e-6;
                              theStep0U2V2: Real from Standard = 1.0e-6)
    returns Boolean from Standard
    is private;
    -- Finds one intersection point of two given surfaces with given 
    --  initial point.
  
  DistanceMinimizeByExtrema(me          : in out;
                            theASurf1   : HSurface from Adaptor3d ;
                            theP0       : Pnt from gp;
                            theU0, theV0: out Real from Standard;
                            theStep0U: Real from Standard = 1.0;
                            theStep0V: Real from Standard = 1.0)
    returns Boolean from Standard
    is private;
    -- Finds one intersection point of two given surfaces with given 
    --  initial point.
  
  SeekPointOnBoundary(me    : in out;
                      theASurf1 , theASurf2  : HSurface from Adaptor3d ;
                      theU1, theV1, theU2, theV2: Real from Standard;
                      isTheFirst : Boolean from Standard)
    returns Boolean from Standard
    is private;
    -- Unites and correctly coordinates of work of
    -- "DistanceMinimizeByGradient" and "DistanceMinimizeByExtrema" functions.
  
  
  PutToBoundary( me    : in out;
                 theASurf1 , theASurf2  : HSurface from Adaptor3d)
    -- Tries to extend existing intersection line 
    --  (as set of points) to surface's boundaries,
    --  if it is possibly.
    --  If line is scienter far from boundaries
    --  or is (almost) parralel with some boundary,
    --  extending is not required.
    returns Boolean from Standard;


  SeekAdditionalPoints( me    : in out;
                        theASurf1 , theASurf2  : HSurface from Adaptor3d;
                        theMinNbPoints : Integer from Standard)
    returns Boolean from Standard;
    -- Unites and correctly coordinates of work of
    -- "DistanceMinimizeByGradient" and "DistanceMinimizeByExtrema" functions.

fields

    done               : Boolean  from Standard;
    line               : LineOn2S from IntSurf;
    close              : Boolean  from Standard;
    tgfirst            : Boolean  from Standard;
    tglast             : Boolean  from Standard;
    indextg            : Integer  from Standard;
    tgdir              : Dir      from gp;

    fleche             : Real     from Standard;   -- max possible vector
    pasMax             : Real     from Standard;   -- max possible uv ratio
    tolconf            : Real     from Standard;   -- tol of confusion of 2 points
    myTolTang          : Real     from Standard;
    pasuv              : Real     from Standard[4];-- uv step on squares 
    pasSav             : Real     from Standard[4];-- first saved step
    pasInit            : Real     from Standard[4];-- saving of steps  
    myStepMin          : Real     from Standard[4];

    Um1                : Real from Standard;
    UM1                : Real from Standard;
    Vm1                : Real from Standard;
    VM1                : Real from Standard;    
    
    Um2                : Real from Standard;
    UM2                : Real from Standard;
    Vm2                : Real from Standard;
    VM2                : Real from Standard;  
    
    ResoU1             : Real from Standard;
    ResoU2             : Real from Standard;
    ResoV1             : Real from Standard;
    ResoV2             : Real from Standard;

    sensCheminement    : Integer  from Standard;
    choixIsoSav        : ConstIsoparametric  from IntImp; 
                       -- save 1st iso choice
    previousPoint      : PntOn2S  from IntSurf;              
                       -- previous intersection point
    previoustg         : Boolean  from Standard;
    previousd          : Dir      from gp;
    previousd1         : Dir2d    from gp;
    previousd2         : Dir2d    from gp;
    firstd1            : Dir2d    from gp;
    firstd2            : Dir2d    from gp;

    myIntersectionOn2S : TheInt2S from IntWalk;
    STATIC_BLOCAGE_SUR_PAS_TROP_GRAND : Integer from Standard;
    STATIC_PRECEDENT_INFLEXION        : Integer from Standard;
end PWalking;
