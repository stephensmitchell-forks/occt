-- Created by: Alexander GRIGORIEV
-- Copyright (c) 2007-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentSection from BinLDrivers

    ---Purpose: More or less independent part of the saved/restored document
    --          that is distinct from OCAF data themselves but may be referred
    --          by them.

uses
    AsciiString      from TCollection,
    Size             from Standard,
    IODevice         from Storage

is
    -- ===== Public methods =====

    Create returns DocumentSection from BinLDrivers;
    ---Purpose: Empty constructor

    Create (theName    : AsciiString from TCollection;
            isPostRead : Boolean from Standard)
        returns DocumentSection from BinLDrivers;
    ---Purpose: Constructor

    Name        (me)
        returns AsciiString from TCollection;
    ---C++: return const&
    ---Purpose: Query the name of the section.

    IsPostRead  (me)
        returns Boolean from Standard;
    ---Purpose: Query the status: if the Section should be read after OCAF;
    --          False means that the Section is read before starting to
    --          read OCAF data.

    Offset      (me)
        returns Size from Standard;
    ---Purpose: Query the offset of the section in the persistent file

    SetOffset   (me:in out; theOffset: Size from Standard);
    ---Purpose: Set the offset of the section in the persistent file

    Length      (me)
        returns Size from Standard;
    ---Purpose: Query the length of the section in the persistent file

    SetLength   (me:in out; theLength: Size from Standard);
    ---Purpose: Set the length of the section in the persistent file

    WriteTOC    (me: in out; theDevice : IODevice from Storage);
    ---Purpose: Create a Section entry in the Document TOC (list of sections)

    Write       (me: in out; theDevice : IODevice from Storage;
                             theOffset: Size from Standard);
    ---Purpose: Save Offset and Length data into the Section entry
    --          in the Document TOC (list of sections)

    ReadTOC     (myclass; theSection: out DocumentSection from BinLDrivers;
                          theDevice : IODevice from Storage);
    ---Purpose: Fill a DocumentSection instance from the data that are read
    --          from TOC.

fields

    myName       : AsciiString from TCollection;
    myValue      : Size from Standard [2];
    myIsPostRead : Boolean from Standard;

end DocumentSection;
