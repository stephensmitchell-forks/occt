-- Created on: 1997-02-06
-- Created by: Kernel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RootData from Storage

inherits TShared from MMgt

uses SequenceOfAsciiString from TColStd,
     AsciiString from TCollection,
     MapOfPers from Storage,
     HSeqOfRoot from Storage,
     Error from Storage,
     Root from Storage
     
raises NoSuchObject from Standard

is

    Create returns RootData from Storage;
    
    NumberOfRoots(me) returns Integer from Standard;
    ---Purpose: returns the number of roots.

    AddRoot(me : mutable;  aRoot : Root from Storage);
    ---Purpose: add a root to <me>. If a root with same name is present, it
    --          will be replaced by <aRoot>.
    
    Roots(me) returns HSeqOfRoot from Storage;
    
    Find(me; aName : AsciiString from TCollection) returns Root from Storage;
    ---Purpose: find a root with name <aName>.
    
    IsRoot(me; aName : AsciiString from TCollection) returns Boolean from Standard;
    ---Purpose: returns Standard_True if <me> contains a root named <aName>
    
    RemoveRoot(me : mutable; aName : AsciiString from TCollection);
    ---Purpose: remove the root named <aName>.

    ErrorStatus(me) returns Error from Storage;
    ErrorStatusExtension(me) returns AsciiString from TCollection;
    
    ClearErrorStatus(me : mutable);
    
    -- PRIVATE

    UpdateRoot(me : mutable; aName : AsciiString from TCollection; aPers : Persistent from Standard) 
    raises NoSuchObject;

    SetErrorStatus(me : mutable; anError : Error from Storage) is private;
    SetErrorStatusExtension(me : mutable; anErrorExt : AsciiString from TCollection) is private;    

    fields
    
      myObjects            : MapOfPers from Storage;
      myErrorStatus        : Error from Storage;
      myErrorStatusExt     : AsciiString      from TCollection;
      
    friends class Schema from Storage
    
end;
