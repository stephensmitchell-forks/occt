-- Created on: 1994-11-30
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeStepWire from TopoDSToStep 
    inherits Root from TopoDSToStep

    ---Purpose: This class implements the mapping between classes 
    --          Wire from TopoDS and TopologicalRepresentationItem from
    --          StepShape. 
  
uses Wire                          from TopoDS,
     TopologicalRepresentationItem from StepShape,
     Tool                          from TopoDSToStep,
     MakeWireError                 from TopoDSToStep,
     FinderProcess_Handle          from Transfer
          
raises NotDone from StdFail
     
is 

    Create returns MakeStepWire;
    
    Create (W : Wire from TopoDS;
    	    T : in out Tool from TopoDSToStep;
	   FP : FinderProcess_Handle from Transfer)
         returns MakeStepWire;
    
    Init(me : in out;
	 W  : Wire from TopoDS;
         T  : in out Tool from TopoDSToStep;
	 FP : FinderProcess_Handle from Transfer);

	    
    Value (me) returns TopologicalRepresentationItem from StepShape
    	raises NotDone
    	is static;
    	---C++: return const&
        
    Error(me) returns MakeWireError from TopoDSToStep;

fields

    myResult : TopologicalRepresentationItem from StepShape;

    myError  : MakeWireError from TopoDSToStep;
    
end MakeStepWire;


