-- Created on: 1996-02-13
-- Created by: Yves FRICAUD
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MakeThickSolid from BRepOffsetAPI inherits MakeOffsetShape from BRepOffsetAPI

	---Purpose: Describes functions to build hollowed solids.
    	-- A hollowed solid is built from an initial solid and a set of
    	-- faces on this solid, which are to be removed. The
    	-- remaining faces of the solid become the walls of the
    	-- hollowed solid, their thickness defined at the time of construction.
    	--        the solid is built from an initial
	--          solid  <S> and a  set of  faces {Fi} from  <S>,
	--          builds a   solid  composed  by two shells closed  by
	--          the {Fi}. First shell <SS>   is composed by all
	--          the faces of <S> expected {Fi}.  Second shell is
	--          the offset shell of <SS>.
    	-- A MakeThickSolid object provides a framework for:
    	-- - defining the cross-section of a hollowed solid,
    	-- - implementing the construction algorithm, and
    	-- - consulting the result.
uses

    MakeOffset  from BRepOffset,
    Mode        from BRepOffset,
    Shape       from TopoDS,
    Face        from TopoDS,
    ListOfShape from TopTools,	
    JoinType    from GeomAbs
    
is


    Create returns MakeThickSolid from BRepOffsetAPI;

    
    Create ( S            : Shape       from TopoDS;
    	     ClosingFaces : ListOfShape from TopTools;
             Offset       : Real        from Standard;
	     Tol          : Real        from Standard  ;
	     Mode         : Mode        from BRepOffset = BRepOffset_Skin;
    	     Intersection : Boolean     from Standard   = Standard_False;
	     SelfInter    : Boolean     from Standard   = Standard_False;
             Join         : JoinType    from GeomAbs    = GeomAbs_Arc;
             RemoveIntEdges : Boolean   from Standard   = Standard_False)
    	---Purpose:  Constructs a hollowed solid from
    	-- the solid S by removing the set of faces ClosingFaces from S, where:
    	--       Offset defines the thickness of the walls. Its sign indicates
    	--   which side of the surface of the solid the hollowed shape is built on;
    	--  - Tol defines the tolerance criterion for coincidence in generated shapes;
    	--  - Mode defines the construction type of parallels applied to free
    	--   edges of shape S. Currently, only one construction type is
    	--   implemented, namely the one where the free edges do not generate
    	--   parallels; this corresponds to the default value BRepOffset_Skin;
    	--   Intersection specifies how the algorithm must work in order to
    	--   limit the parallels to two adjacent shapes:
    	-- - if Intersection is false (default value), the intersection
    	--   is calculated with the parallels to the two adjacent shapes,
    	--  -     if Intersection is true, the intersection is calculated by
    	--   taking account of all parallels generated; this computation
    	--   method is more general as it avoids self-intersections
    	--   generated in the offset shape from features of small dimensions
    	--   on shape S, however this method has not been completely
    	--   implemented and therefore is not recommended for use;
    	--  -     SelfInter tells the algorithm whether a computation to
    	--   eliminate self-intersections needs to be applied to the
    	--   resulting shape. However, as this functionality is not yet
    	--   implemented, you should use the default value (false);
    	--  - Join defines how to fill the holes that may appear between
    	--   parallels to the two adjacent faces. It may take values
    	--   GeomAbs_Arc or GeomAbs_Intersection:
    	-- - if Join is equal to GeomAbs_Arc, then pipes are generated
    	--           between two free edges of two adjacent parallels,
    	--           and spheres are generated on "images" of vertices;
    	--           it is the default value,
    	-- - if Join is equal to GeomAbs_Intersection,
    	--   then the parallels to the two adjacent faces are
    	--   enlarged and intersected, so that there are no free
    	--   edges on parallels to faces.
    	--   Warnings
    	-- Since the algorithm of MakeThickSolid is based on
    	-- MakeOffsetShape algorithm, the warnings are the same as for
    	-- MakeOffsetShape.
    returns MakeThickSolid from BRepOffsetAPI;
    
    Build (me : in out)
    is redefined;
	---Purpose: Builds the resulting shape (redefined from MakeOffsetShape).
	---Level: Public     


    Modified (me: in out; S : Shape from TopoDS)
    	---Purpose: Returns the list  of shapes modified from the shape
    	--          <S>. 
        ---C++: return const & 
        ---Level: Public
    returns ListOfShape from TopTools
    is redefined virtual;


end MakeThickSolid;
