-- Created by: Peter KURNEV
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

class BOP from BOPAlgo  
    inherits Builder from BOPAlgo
---Purpose: 

uses
    Shape from TopoDS,  
    BaseAllocator from BOPCol,  
    ListOfShape from BOPCol, 
    MapOfShape  from BOPCol,  
    --modified by NIZHNY-EMV Fri Sep 02 08:38:28 2011 
    IndexedDataMapOfShapeListOfShape from BOPCol,
    --modified by NIZHNY-EMV Fri Sep 02 08:38:30 2011 
    Operation from BOPAlgo, 
    PaveFiller from BOPAlgo 

--raises

is
    Create 
    ---Purpose:  Empty constructor     
    returns BOP from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_BOP();"  
      
    Create (theAllocator: BaseAllocator from BOPCol)
    returns BOP from BOPAlgo; 
	 
    Clear(me:out) 
    is redefined; 
    ---Purpose:  Clears internal fields and arguments   
     
    AddArgument (me:out;  
        theShape: Shape from TopoDS) 
    ---Purpose:  Adds Object argument of the operation     
     is redefined;
	 
    AddTool (me:out;  
        theShape: Shape from TopoDS) 
    ---Purpose:  Adds Tool argument of the operation    	     
    is virtual; 
	 
    Object(me) 
    returns Shape from TopoDS; 
    ---C++: return const &   

    Tool(me) 
    returns Shape from TopoDS; 
    ---C++: return const &   

    SetOperation(me:out;  
        theOperation: Operation from BOPAlgo); 
	 
    Operation(me) 
    returns Operation from BOPAlgo;  
    --
    --  protected methods 
    -- 
    CheckData(me:out) 
    is redefined protected; 

    Prepare(me:out)  
    is redefined protected; 
    ---Purpose:  Provides preparing actions 

    PerformInternal(me:out; 
        thePF:PaveFiller from BOPAlgo) 
    is redefined protected;   
    ---Purpose:  Performs calculations using prepared Filler 
    --           object theDSF          	 
      
    BuildShape(me:out) 
    is protected; 
 
    BuildRC(me:out) 
    is protected; 
 
    BuildSolid(me:out) 
    is protected; 
	 
    BuildSection(me:out) 
    is protected;  
     
    Dimension(myclass; 
        theS:Shape from TopoDS) 
    returns Integer from Standard;
    --is protected;  
	 
    TreatCompound(myclass; 
        theS:Shape from TopoDS; 
        theLS:out ListOfShape from BOPCol) 
    is protected;     
     
    --modified by NIZHNY-EMV Fri Sep 02 08:34:17 2011 
    IsBoundSplits(me:out; 
        theS:Shape from TopoDS; 
        theMEF:out IndexedDataMapOfShapeListOfShape from BOPCol)  
    returns Boolean from Standard
    is protected;
    --modified by NIZHNY-EMV Fri Sep 02 08:34:19 2011

fields 
    myNbArgs    : Integer from Standard    is protected;
    myOperation : Operation from BOPAlgo   is protected; 
    myArgs      : Shape from TopoDS[2]     is protected;  
    myDims      : Integer from Standard[2] is protected;  
    -- 
    myRC        : Shape from TopoDS        is protected; 
    myTools     : ListOfShape from BOPCol  is protected; 
    myMapTools  : MapOfShape  from BOPCol  is protected;  
    
end BOP;
