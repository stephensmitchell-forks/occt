-- Created on: 2000-08-16
-- Created by: Andrey BETENEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IGESCAFControl 

    ---Purpose: Provides high-level API to translate IGES file
    --          to and from DECAF document

uses
    Quantity,
    TCollection,
    TopoDS,
    TopTools,
    TDocStd,
    TDF,
    XCAFDoc,
    XCAFPrs,
    XSControl,
    IGESControl

is

    imported Reader;
    	---Purpose: Provides a tool for reading IGES file

    imported Writer;
    	---Purpose: Provides a tool for writing IGES file

    DecodeColor (col: Integer) returns Color from Quantity;
    	---Purpose: Converts IGES color index to CASCADE color

    EncodeColor (col: Color from Quantity) returns Integer;
    	---Purpose: Tries to Convert CASCADE color to IGES color index
	--          If no corresponding color defined in IGES, returns 0
	

end IGESCAFControl;
