-- Created on: 1995-03-06
-- Created by: Laurent PAINNOT
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package Poly

        ---Purpose: This  package  provides  classes  and services  to
        --          handle :
        --
        --          * 3D triangular polyhedrons.
        --
        --          * 3D polygons.
        --
        --          * 2D polygon.
        --
        --          * Tools to dump, save and restore those objects.

uses

    MMgt,
    TCollection,
    TColStd,
    gp,
    TColgp,
    TShort

is

    class Triangle;

    class Array1OfTriangle
    instantiates Array1 from TCollection(Triangle from Poly);

    class HArray1OfTriangle
    instantiates HArray1 from TCollection(Triangle         from Poly,
                                          Array1OfTriangle from Poly);

    imported transient class Triangulation;
    imported transient class Mesh;
    imported Element;

    class Polygon3D;

    class Polygon2D;

    class PolygonOnTriangulation;

    --
    -- Tools to use triangulations
    --

    class Connect;
        ---Purpose: Computes and  stores  the    link from   nodes  to
        --          triangles     and from triangles to   neighbouring
        --          triangles.
        -- This tool is obsolete, replaced by Poly_CoherentTriangulation

    --
    --     Data types for the Coherent Triangulation data model
    --
    imported CogerentTriangulation;
    imported CoherentTriangle;
    imported CoherentNode;
    imported CoherentLink;
    imported CoherentTriPtr;
    imported ListOfTriangulation;

    imported MakeLoops;
        ---Purpose: Algorithm to make minimal loops in a graph

    --
    --  Package methods
    --

    Catenate (lstTri: ListOfTriangulation from Poly)
        returns Triangulation from Poly;
        ---Purpose: Join several triangulations to one new triangulation object.
        --          The new triangulation is just a mechanical sum of input
        --          triangulations, without node sharing. UV coordinates are
        --          dropped in the result.

    Write(T       : Triangulation from Poly;
          OS      : in out OStream;
          Compact : Boolean = Standard_True);

        ---Purpose: Writes the content of the triangulation <T> on the
        --          stream <OS>. If <Compact> is true this is a "save"
        --          format  intended  to  be read back   with the Read
        --          method. If compact is False  it is a "Dump" format
        --          intended to be informative.

    Write(P       : Polygon3D from Poly;
          OS      : in out OStream;
          Compact : Boolean = Standard_True);

        ---Purpose: Writes  the  content  of the 3D polygon <P> on the
        --          stream <OS>. If <Compact> is true this is a "save"
        --          format  intended  to  be read back   with the Read
        --          method. If compact is False  it is a "Dump" format
        --          intended to be informative.

    Write(P       : Polygon2D from Poly;
          OS      : in out OStream;
          Compact : Boolean = Standard_True);

        ---Purpose: Writes the  content  of the 2D polygon  <P> on the
        --          stream <OS>. If <Compact> is true this is a "save"
        --          format  intended  to  be read back   with the Read
        --          method. If compact is False  it is a "Dump" format
        --          intended to be informative.


    Dump(T       : Triangulation from Poly;
         OS      : in out OStream);
       ---Purpose: Dumps  the triangulation.  This   is a call to  the
       --          previous method with Comapct set to False.

    Dump(P       : Polygon3D from Poly;
         OS      : in out OStream);
       ---Purpose: Dumps  the  3D  polygon.  This   is a call to  the
       --          previous method with Comapct set to False.

    Dump(P       : Polygon2D from Poly;
         OS      : in out OStream);
       ---Purpose: Dumps  the  2D  polygon.  This   is a call to  the
       --          previous method with Comapct set to False.


    ReadTriangulation(IS : in out IStream)
    returns Triangulation from Poly;
        ---Purpose: Reads a triangulation from the stream <IS>.

    ReadPolygon3D(IS : in out IStream)
    returns Polygon3D from Poly;
        ---Purpose: Reads a 3d polygon from the stream <IS>.

    ReadPolygon2D(IS : in out IStream)
    returns Polygon2D from Poly;
        ---Purpose: Reads a 2D polygon from the stream <IS>.

    ComputeNormals(Tri : Triangulation from Poly);
        ---Purpose: Compute node normals for face triangulation
        --  as mean normal of surrounding triangles

    PointOnTriangle(P1, P2, P3, P: XY from gp; UV: out XY from gp)
    returns Real;
        ---Purpose: Computes parameters of the point P on triangle
        --          defined by points P1, P2, and P3, in 2d.
        --          The parameters U and V are defined so that
        --          P = P1 + U * (P2 - P1) + V * (P3 - P1),
        --          with U >= 0, V >= 0, U + V <= 1.
        --          If P is located outside of triangle, or triangle
        --          is degenerated, the returned parameters correspond
        --          to closest point, and returned value is square of
        --          the distance from original point to triangle (0 if
        --          point is inside).

end Poly;
