-- Created on: 2004-01-09
-- Created by: Sergey KUUL
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Dimension from XCAFDoc inherits Attribute from TDF

	---Purpose: attribute to store dimension

uses
    Label from TDF,
    RelocationTable from TDF,
    DimensionObject from XCAFDimTolObjects

is

    Create returns Dimension from XCAFDoc;
    
    ---Category: class methods
    --           =============

    GetID (myclass)   
    	---C++: return const &  
    returns GUID from Standard;
    
    Set (myclass; theLabel : Label from TDF)
    returns Dimension from XCAFDoc;
                                                                          
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; With : Attribute from TDF);

    NewEmpty (me)
    returns Attribute from TDF;

    Paste (me; Into : Attribute from TDF;
	       RT   : RelocationTable from TDF);    

    SetObject (me : mutable; theDimensionObject : DimensionObject from XCAFDimTolObjects);

    GetObject (me) returns DimensionObject from XCAFDimTolObjects;

end Dimension;
