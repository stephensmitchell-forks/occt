-- Created by: Peter KURNEV
-- Copyright (c) 2010-2012 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class FaceInfo from BOPDS 

	---Purpose: 
    	-- The class BOPDS_FaceInfo is to store  
    	-- handy information about state of face
uses     
    BaseAllocator from BOPCol,
    MapOfInteger from BOPCol,
    MapOfPaveBlock from BOPDS
   
--raises

is
    Create 
    	returns FaceInfo from BOPDS; 
    ---C++: inline 	 
    ---C++: alias "virtual ~BOPDS_FaceInfo();"  
      	---Purpose:  
    	--- Empty contructor  
    	---   
	 
    Create (theAllocator: BaseAllocator from BOPCol) 
    	returns FaceInfo from BOPDS;  
    ---C++: inline   
    	---Purpose:   
     	---  Contructor    
    	---  theAllocator - the allocator to manage the memory     
    	---    
	
    Clear(me:out); 
    	---Purpose:   
     	---  Clears the contents      
    
    SetIndex(me:out; 
    	    theI: Integer from Standard); 
    ---C++: inline 
     	---Purpose: 
    	--- Modifier   
	--- Sets the index of the face <theI> 
	
    Index(me) 
    	returns Integer from Standard; 
    ---C++: inline  
    	---Purpose: 
    	--- Selector   
	--- Returns the index of the face 
    --  
    -- In 
    --  
    PaveBlocksIn(me) 
	returns MapOfPaveBlock from BOPDS; 
    ---C++: return const &  
    ---C++: inline 
     	---Purpose: 
    	--- Selector   
	--- Returns the pave blocks of the face 
	--- that  have state In 
	 
    ChangePaveBlocksIn(me:out) 
    	returns MapOfPaveBlock from BOPDS;  
    ---C++: return &  
    ---C++: inline    
      	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the pave blocks  
    	--  of the face 
	--- that  have state In 
	 
    VerticesIn(me) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return const &  
    ---C++: inline  
     	---Purpose: 
    	--- Selector   
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state In  
	
    ChangeVerticesIn(me:out) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return &  
    ---C++: inline 
    	---Purpose: 
    	--- Selector/Modifier    
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state In   
    --  
    -- On 
    --  
    PaveBlocksOn(me) 
	returns MapOfPaveBlock from BOPDS; 
    ---C++: return const &  
    ---C++: inline    
    	---Purpose: 
    	--- Selector   
	--- Returns the pave blocks of the face 
	--- that  have state On
     
    ChangePaveBlocksOn(me:out) 
    	returns MapOfPaveBlock from BOPDS;  
    ---C++: return &  
    ---C++: inline    
      	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the pave blocks  
    	--  of the face 
	--- that  have state On 
    VerticesOn(me) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return const &  
    ---C++: inline  
     	---Purpose: 
    	--- Selector   
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state On 
	 
    ChangeVerticesOn(me:out) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return &  
    ---C++: inline 
    	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the list of indices for vertices  
    	--  of the face
	--- that have state On   
    --  
    -- Sections 
    --  
    PaveBlocksSc(me) 
	returns MapOfPaveBlock from BOPDS; 
    ---C++: return const &  
    ---C++: inline   
    	---Purpose: 
    	--- Selector   
	--- Returns the pave blocks of the face 
	--- that are  pave blocks of section edges  
     
    ChangePaveBlocksSc(me:out) 
    	returns MapOfPaveBlock from BOPDS;  
    ---C++: return &  
    ---C++: inline  
    	--- Selector/Modifier      
	--- Returns the pave blocks of the face 
	--- that are  pave blocks of section edges     
      
    VerticesSc(me) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return const &  
    ---C++: inline  
    	---Purpose: 
    	--- Selector   
	--- Returns the list of indices for section  vertices  
    	--  of the face
     
    ChangeVerticesSc(me:out) 
    	returns MapOfInteger from BOPCol;  
    ---C++: return &  
    ---C++: inline 
    	---Purpose: 
    	--- Selector/Modifier   
	--- Returns the list of indices for section  vertices  
    	--  of the face 
    --  
    -- Others
    --    
    --Update(me:out) 
    --	is protected; 
     
fields 
    myAllocator   : BaseAllocator from BOPCol is protected; 
    myIndex       : Integer from Standard is protected; 
    myPaveBlocksIn: MapOfPaveBlock from BOPDS is protected;  
    myVerticesIn  : MapOfInteger from BOPCol is protected;  
    myPaveBlocksOn: MapOfPaveBlock from BOPDS is protected;  
    myVerticesOn  : MapOfInteger from BOPCol is protected;
    myPaveBlocksSc: MapOfPaveBlock from BOPDS is protected;  
    myVerticesSc  : MapOfInteger from BOPCol is protected;
 
end FaceInfo;
