-- Created by: Peter KURNEV
-- Copyright (c) 2010-2014 OPEN CASCADE SAS
-- Copyright (c) 2007-2010 CEA/DEN, EDF R&D, OPEN CASCADE
-- Copyright (c) 2003-2007 OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN, CEDRAT,
--                         EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PaveFiller from BOPAlgo 
   inherits Algo from BOPAlgo 
    ---Purpose: 

uses 
    Pnt from gp,  
    ShapeEnum from TopAbs,  
    Vertex from TopoDS,
    Face from TopoDS, 
    Edge from TopoDS,  
        
    ListOfShape from TopTools,
     
    BaseAllocator from BOPCol, 
    ListOfShape from BOPCol, 
    MapOfInteger from BOPCol, 
    ListOfInteger from BOPCol, 
    DataMapOfShapeInteger from BOPCol,   
    IndexedDataMapOfShapeInteger from BOPCol,   
    DataMapOfIntegerListOfInteger from BOPCol, 
    DataMapOfShapeListOfShape from BOPCol,
    IndexedDataMapOfShapeListOfShape from BOPCol, 
    DataMapOfIntegerReal from BOPCol, 
    DataMapOfIntegerInteger from BOPCol,
    --  
    Context from IntTools,
    -- 
    SectionAttribute from BOPAlgo, 
    
    DS  from BOPDS,
    PDS from BOPDS, 
    Iterator  from BOPDS, 
    PIterator from BOPDS, 
    PaveBlock from BOPDS, 
    Curve from BOPDS,  
    IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS,
    MapOfPaveBlock from BOPDS,  
    IndexedMapOfPaveBlock from BOPDS,  
    ListOfPaveBlock from BOPDS, 
    ListOfPave from BOPDS, 
    ListOfPntOn2S from IntSurf, 
    Curve from IntTools,
    
    DataMapOfPaveBlockListOfPaveBlock from BOPDS, 
    VectorOfCurve from BOPDS 
     
--raises

is 
    Create 
      returns PaveFiller from BOPAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~BOPAlgo_PaveFiller();"
     
    Create (theAllocator: BaseAllocator from BOPCol) 
      returns PaveFiller from BOPAlgo;   
 
    DS(me:out) 
      returns DS from BOPDS; 
    ---C++:return  const &   
    
      
    PDS(me:out) 
      returns PDS from BOPDS; 
     
    Iterator(me:out) 
      returns PIterator from BOPDS;  
    ---C++:return const & 
     
    SetArguments(me:out; 
            theLS:ListOfShape from BOPCol);   
            
    SetArguments(me:out; 
            theLS:ListOfShape from TopTools);  

    Arguments(me) 
      returns ListOfShape from BOPCol; 
    ---C++: return const & 

    Context(me:out) 
      returns Context from IntTools;  
       
    SetSectionAttribute(me:out; 
        theSecAttr : SectionAttribute from BOPAlgo); 
         
    Perform(me:out) 
      is redefined;   
    --  
    -- protected methods 
    --  
    PerformInternal (me:out) 
      is virtual protected;   
      
    Clear(me:out) 
      is virtual protected;  
          
    Init(me:out) 
      is virtual protected;
     
    Prepare(me:out) 
      is  protected;
     
    PerformVV(me:out) 
      is virtual protected;   
     
    PerformVE(me:out) 
      is virtual protected;  
     
    PerformVF(me:out) 
      is virtual protected;  
  
    PerformEE(me:out) 
      is virtual protected; 
   
    PerformEF(me:out) 
      is virtual protected; 
     
    PerformFF(me:out) 
      is virtual protected;
     
    PerformVZ(me:out) 
      is virtual protected; 
       --Purpose: Computes Vertex/Solid interferences 
       
    PerformEZ(me:out) 
      is virtual protected;  
      --Purpose: Computes Edge/Solid interferences 
     
    PerformFZ(me:out) 
      is virtual protected;   
      --Purpose: Computes Face/Solid interferences 
    PerformZZ(me:out) 
      is virtual protected;  
      --Purpose: Computes Solid/Solid interferences  
  
    PerformSZ(me:out; 
        aTS:ShapeEnum from TopAbs) 
      is virtual protected;
 
    TreatVerticesEE(me:out) 
      is protected; 

    MakeSplitEdges(me:out) 
      is protected;   
        
    MakeBlocks(me:out) 
      is protected; 
  
    MakePCurves(me:out) 
      is protected; 
  
    ProcessDE(me:out) 
      is protected;  
       
    FillShrunkData(me:out; 
        thePB:out PaveBlock from BOPDS) 
      is protected;   
 
    FillShrunkData(me:out; 
        theType1: ShapeEnum from TopAbs; 
        theType2: ShapeEnum from TopAbs) 
      is protected;   
 
    PerformVerticesEE(me:out; 
        theMVCPB:out IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol) 
      returns Integer from Standard 
      is protected; 
  
    PerformVerticesEF(me:out; 
        theMVCPB:out IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS; 
        theAllocator:out BaseAllocator from BOPCol) 
      returns Integer from Standard 
      is protected; 
     
    CheckFacePaves(me:out; 
        theVnew:Vertex from TopoDS; 
        theMIF:MapOfInteger from BOPCol) 
      returns Boolean from Standard 
      is protected;  
   
    CheckFacePaves(myclass; 
        theN:Integer from Standard; 
        theMIFOn:MapOfInteger from BOPCol; 
        theMIFIn:MapOfInteger from BOPCol) 
      returns Boolean from Standard 
      is protected;  
  
    IsExistingVertex(me; 
        theP:Pnt from gp; 
        theTol:Real from Standard; 
        theMVOn:MapOfInteger from BOPCol) 
      returns Boolean from Standard 
      is protected; 

    PutPavesOnCurve(me:out; 
        theMVOn   : MapOfInteger from BOPCol; 
        theTolR3D : Real from Standard; 
        theNC     : out Curve from BOPDS;  
        nF1       : Integer from Standard; 
        nF2       : Integer from Standard; 
        theMI     : MapOfInteger from BOPCol; 
        theMVEF   : MapOfInteger from BOPCol; 
        theMVTol  : out DataMapOfIntegerReal from BOPCol) 
      is protected;   
    ---Purpose: 
    -- Checks and puts paves from <theMVOn> on the curve <theNC>.

    ExtendedTolerance(me:out; 
        nV       : Integer from Standard; 
        aMI      : MapOfInteger from BOPCol; 
        aTolVExt : out Real from  Standard;
        aType    : Integer from Standard = 0) 
      returns Boolean from  Standard 
      is protected; 
    ---Purpose: 
    -- Depending on the parameter aType it checks whether  
    -- the vertex nV was created in EE or EF intersections. 
    -- If so, it increases aTolVExt from tolerance value of vertex to  
    -- the max distance from vertex nV to the ends of the range of common part. 
    -- Possible values of aType: 
    -- 1 - checks only EE; 
    -- 2 - checks only EF;
    -- other - checks both types of intersections.
  
    PutBoundPaveOnCurve(me:out;  
        theF1: Face from TopoDS;  
        theF2: Face from TopoDS;  
        theTolR3D:Real from Standard; 
        theNC:out Curve from BOPDS;  
        theLBV:out ListOfInteger from BOPCol) 
      is protected; 

    IsExistingPaveBlock(me:out; 
        thePB:PaveBlock from BOPDS;  
        theNC:Curve from BOPDS;
        theTolR3D:Real from Standard; 
        theMPB:IndexedMapOfPaveBlock from BOPDS; 
        thePBOut:out PaveBlock from BOPDS)
      returns Boolean from Standard 
      is protected;  
 
    IsExistingPaveBlock(me:out; 
        thePB:PaveBlock from BOPDS;  
        theNC:Curve from BOPDS;
        theLSE:ListOfInteger from BOPCol) 
      returns Boolean from Standard 
      is protected;   
     
    PostTreatFF(me:out; 
        theMSCPB:out IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS; 
        theMVI:out DataMapOfShapeInteger from BOPCol;  
        theDMExEdges:out DataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theDMI:out DataMapOfIntegerInteger from BOPCol;
        theAllocator:out BaseAllocator from BOPCol) 
      returns Integer from Standard 
      is protected;  
    ---Purpose: 
    -- Treatment of section edges.
    
    --
    --  Treatment of degenerated edges  
    -- 
    FindPaveBlocks(me:out;  
        theV:Integer from Standard; 
        theF:Integer from Standard; 
        theLPB:out ListOfPaveBlock from BOPDS) 
      is protected; 

    FillPaves(me:out;  
        theV:Integer from Standard; 
        theE:Integer from Standard; 
        theF:Integer from Standard; 
        theLPB: ListOfPaveBlock from BOPDS; 
        thePB: PaveBlock from BOPDS) 
      is protected; 
  
    MakeSplitEdge(me:out;  
        theV:Integer from Standard; 
        theF:Integer from Standard) 
      is protected;  
      
    GetEFPnts(me:out;
        nF1 : Integer from Standard;
        nF2 : Integer from Standard;
        aListOfPnts: out ListOfPntOn2S from IntSurf)
      is protected; 
       
    PutEFPavesOnCurve(me:out; 
        theNC      : out Curve from BOPDS; 
        theMI      : MapOfInteger from BOPCol;
        theMVEF    : MapOfInteger from BOPCol;
        theMVTol   : out DataMapOfIntegerReal from BOPCol)
      is protected; 
    ---Purpose: 
    -- Checks and puts paves created in EF intersections on the curve <theNC>.
 
    PutStickPavesOnCurve(me:out; 
        aF1        : Face from TopoDS; 
        aF2        : Face from TopoDS;  
        theMI      : MapOfInteger from BOPCol;
        theNC      : out Curve from BOPDS; 
        theMVStick : MapOfInteger from BOPCol; 
        theMVTol   : out DataMapOfIntegerReal from BOPCol)
      is protected;  
    ---Purpose: 
    -- Puts stick paves on the curve <theNC>
 
    GetStickVertices(me:out; 
        nF1        : Integer from Standard; 
        nF2        : Integer from Standard; 
        theMVStick : out MapOfInteger from BOPCol;
        theMVEF    : out MapOfInteger from BOPCol; 
        theMI      : out MapOfInteger from BOPCol)
      is protected;  
    ---Purpose: 
    -- Collects indices of vertices created in all intersections between 
    -- two faces (<nF1> and <nF2>) to the map <theMVStick>. 
    -- Also, it collects indices of EF vertices to the <theMVEF> map  
    -- and indices of all subshapes of these two faces to the <theMI> map.
 
    GetFullShapeMap(me:out; 
        nF    : Integer from Standard; 
        theMI : out MapOfInteger from BOPCol) 
      is protected; 
    ---Purpose: 
    -- Collects index nF and indices of all subshapes of the shape with index <nF>
    -- to the map <theMI>. 
    
    RemoveUsedVertices(me:out; 
        theNC : out Curve from BOPDS; 
        theMV : out MapOfInteger from BOPCol)  
      is protected; 
    ---Purpose: 
    -- Removes indices of vertices that are already on the
    -- curve <theNC> from the map <theMV>.  
    -- It is used in PutEFPavesOnCurve and PutStickPavesOnCurve methods.
 
    PutPaveOnCurve(me:out; 
        nV        : Integer from Standard; 
        theTolR3D : Real from Standard;
        theNC     : out Curve from BOPDS; 
        theMI     : MapOfInteger from BOPCol;
        theMVTol  : out DataMapOfIntegerReal from BOPCol;
        aType     : Integer from Standard = 0)
      is protected; 
    ---Purpose: 
    -- Puts the pave nV on the curve theNC.  
    -- Parameter aType defines whether to check the pave with 
    -- extended tolerance: 
    -- 0 - do not perform the check; 
    -- other - perform the check (aType goes to ExtendedTolerance).
 
    ProcessExistingPaveBlocks(me:out; 
        theInt     : Integer from Standard; 
        theMPBOnIn : IndexedMapOfPaveBlock from BOPDS; 
        theDMBV    : DataMapOfIntegerListOfInteger from BOPCol; 
        theMSCPB   : out IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS; 
        theMVI     : out DataMapOfShapeInteger from BOPCol; 
        theMPB     : out MapOfPaveBlock from BOPDS)
      is  protected; 
    ---Purpose:       
    -- Adds the existing edges from the map <theMPBOnIn> which interfere  
    -- with the vertices from <theMVB> map to the post treatment of section edges.
 
    UpdateExistingPaveBlocks(me:out; 
        thePB   : PaveBlock from BOPDS;
        theLPB  : out ListOfPaveBlock from BOPDS; 
        nF1     : Integer from Standard; 
        nF2     : Integer from Standard)
      is protected; 
    ---Purpose: 
    -- Replaces existing pave block <thePB> with new pave blocks <theLPB>. 
    -- The list <theLPB> contains images of <thePB> which were created in 
    -- the post treatment of section edges.
 
    TreatNewVertices(me:out; 
        theMVI    : IndexedDataMapOfShapeInteger from BOPCol; 
        theImages : out IndexedDataMapOfShapeListOfShape from BOPCol) 
      is protected; 
    ---Purpose: 
    -- Treatment of vertices that were created in EE intersections. 
 
    PutClosingPaveOnCurve (me:out; 
        aNC :out Curve from BOPDS)  
      is protected; 
    ---Purpose: 
    -- Put paves on the curve <aBC> in case when <aBC>   
    -- is closed 3D-curve  
     
    PreparePostTreatFF(me:out; 
        aInt   : Integer from Standard;
        aCur   : Integer from Standard;
        aPB    : PaveBlock from BOPDS;  
        aMSCPB : out IndexedDataMapOfShapeCoupleOfPaveBlocks from BOPDS; 
        aMVI   : out DataMapOfShapeInteger from BOPCol; 
        aLPB   : out ListOfPaveBlock from BOPDS)
      is protected; 
    ---Purpose: 
    -- Keeps data for post treatment 
     
    RefineFaceInfoOn(me:out) 
      is protected; 
    ---Purpose: 
    -- Refines the state On for the all faces having 
    -- state information 

    UpdateFaceInfo(me:out;
        theDME:out DataMapOfPaveBlockListOfPaveBlock from BOPDS; 
        theDMV: DataMapOfIntegerInteger from BOPCol) 
      is protected; 
    ---Purpose: 
    -- Updates the information about faces
     
    ForceInterfVE(me:out; 
        nV   : Integer from Standard; 
        aPB  : out PaveBlock from BOPDS; 
        aMPB : out MapOfPaveBlock from BOPDS) 
      is protected;
    ---Purpose: 
    -- Updates tolerance of vertex with index <nV>  
    -- to make it interfere with edge
    
    ForceInterfVF(me:out; 
        nV : Integer from Standard; 
        nF : Integer from Standard) 
      returns Boolean from Standard
      is protected;
    ---Purpose: 
    -- Updates tolerance of vertex with index <nV>  
    -- to make it interfere with face with index <nF> 
    
    CheckPlanes(me; 
        nF1 : Integer from Standard; 
        nF2 : Integer from Standard)
      returns Boolean from Standard 
      is protected; 
    ---Purpose: 
    -- Checks if there are any common or intersecting sub shapes
    -- between two planar faces.  
     
    SplitEdge(me:out; 
        nE  : Integer from Standard; 
        nV1 : Integer from Standard; 
        aT1 : Real from Standard;
        nV2 : Integer from Standard; 
        aT2 : Real from Standard) 
    returns Integer from Standard 
    is protected;
    ---Purpose: 
    -- Creates new edge from the edge nE with vertices nV1 and nV2 
    -- and returns the index of that new edge in the DS.
 
    UpdatePaveBlocks(me:out;  
        theDMI : DataMapOfIntegerInteger from BOPCol) 
    is protected; 
    ---Purpose: 
    -- Updates pave blocks which have the paves with indices contained  
    -- in the map <theDMI>.

    SetFuzzyValue(me:out; 
        theFuzz : Real from Standard);
    ---Purpose: Sets the additional tolerance

    FuzzyValue(me)
    returns Real from Standard;
    ---Purpose: Returns the additional tolerance 

fields  
    myArguments   : ListOfShape from BOPCol is protected;  
    myDS          : PDS from BOPDS is protected; 
    myIterator    : PIterator from BOPDS is protected; 
    myContext     : Context from IntTools is protected;   
    mySectionAttribute : SectionAttribute from BOPAlgo is protected;
    myFuzzyValue  : Real from Standard is protected;
end PaveFiller;
