-- Created on: 1995-06-06
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BRepApprox 

	---Purpose: This package provides services on intersection curves
	--          dealt by topological operations on BRep objects.
	--          Services are approximation services.


uses

    MMgt,
    TColStd,
    gp,
    GeomAbs,
    Adaptor3d,
    Geom,
    Geom2d,
    BRepAdaptor,
    IntSurf,
    ApproxInt
    
is

    class ApproxLine;
	
    class SurfaceTool;
    
    imported Approx;

end BRepApprox;
