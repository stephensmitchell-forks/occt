-- Created on: 2002-12-06
-- Created by: data exchange team
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Construct from StepAP209 inherits Tool from STEPConstruct

    ---Purpose: Basic tool for working with AP209 model

uses
    WorkSession_Handle from XSControl,
    Product from StepBasic,
    ProductDefinition from StepBasic,
    ProductDefinitionFormation from StepBasic,
    ProductDefinitionShape from StepRepr,
    HSequenceOfElementRepresentation from StepFEA,
    HSequenceOfElementMaterial from StepElement,
    HSequenceOfCurveElementSectionDefinition from StepElement,
    HSequenceOfElementGeometricRelationship from StepFEA,
    FeaModel from StepFEA,
    ShapeRepresentation from StepShape,
    Curve3dElementRepresentation from StepFEA,
    ElementRepresentation from StepFEA,
    FeaAxis2Placement3d from StepFEA,
    StepModel from StepData


is

    Create returns Construct;
    	---Purpose: Creates an empty tool

    Create (WS: WorkSession_Handle from XSControl) returns Construct;
    	---Purpose: Creates a tool and initializes it
	
    Init (me: in out; WS: WorkSession_Handle from XSControl) returns Boolean;
    	---Purpose: Initializes tool; returns True if succeeded

    IsDesing(me; PD: ProductDefinitionFormation from StepBasic) returns Boolean;
    IsAnalys(me; PD: ProductDefinitionFormation from StepBasic) returns Boolean;


    -- methods for getting fea_model
    FeaModel(me; Prod: Product from StepBasic) returns FeaModel from StepFEA;

    FeaModel(me; PDF: ProductDefinitionFormation from StepBasic) returns FeaModel from StepFEA;


    -- methods for gettig fea_axis2_placement_3d
    GetFeaAxis2Placement3d(me; theFeaModel: FeaModel from StepFEA)
    returns FeaAxis2Placement3d from StepFEA;


    -- methods for getting idealized_analysis_shape
    IdealShape(me; Prod: Product from StepBasic) returns ShapeRepresentation from StepShape;

    IdealShape(me; PDF: ProductDefinitionFormation from StepBasic) returns ShapeRepresentation from StepShape;


    -- methods for getting nominal_design_shape
    NominShape(me; Prod: Product from StepBasic) returns ShapeRepresentation from StepShape;

    NominShape(me; PDF: ProductDefinitionFormation from StepBasic) returns ShapeRepresentation from StepShape;


    -- method for getting list of element_material
    GetElementMaterial(me) returns HSequenceOfElementMaterial from StepElement;
    
    -- method for getting list of element_geometric_relationship
    GetElemGeomRelat(me) returns HSequenceOfElementGeometricRelationship from StepFEA;
    

    -- methods for getting list of element_representations
    GetElements1D(me; theFeaModel: FeaModel from StepFEA)
    returns HSequenceOfElementRepresentation from StepFEA;
    
    GetElements2D(me; theFEAModel: FeaModel from StepFEA)
    returns HSequenceOfElementRepresentation from StepFEA;
    
    GetElements3D(me; theFEAModel: FeaModel from StepFEA)
    returns HSequenceOfElementRepresentation from StepFEA;

    GetFeaElements(me; theFeaModel: FeaModel from StepFEA;
    	    	       theType: Type from Standard)
    returns HSequenceOfElementRepresentation from StepFEA is protected;


    GetCurElemSection(me; ElemRepr: Curve3dElementRepresentation from StepFEA)
    returns HSequenceOfCurveElementSectionDefinition from StepElement;
    --- Purpose: Getting list of curve_element_section_definitions
    ---          for given element_representation 

    GetShReprForElem(me; ElemRepr: ElementRepresentation from StepFEA)
    returns ShapeRepresentation from StepShape;
        
    CreateAnalysStructure(me; Prod: Product from StepBasic) returns Boolean from Standard;
    --- Purpose: Create empty structure for idealized_analysis_shape

    CreateFeaStructure(me; Prod: Product from StepBasic) returns Boolean from Standard;
    --- Purpose: Create fea structure 

    ReplaceCcDesingToApplied(me) returns Boolean from Standard;
    --- Purpose: Put into model entities Applied... for AP209 instead of
    --           entities CcDesing... from AP203.

    CreateAddingEntities(me; AnaPD: ProductDefinition from StepBasic) returns Boolean from Standard;
    --- Purpose: Create approval.. , date.. , time.. , person.. and
    --           organization.. entities for analysis structure

    CreateAP203Structure(me) returns StepModel from StepData;
    --- Purpose: Create AP203 structure from existing AP209 structure

    CreateAdding203Entities(me; PD: ProductDefinition from StepBasic;
                                aModel: in out StepModel from StepData)
    returns Boolean from Standard;
    --- Purpose: Create approval.. , date.. , time.. , person.. and
    --           organization.. entities for 203 structure

    -- auxiliary methods
    FeaModel(me; PDS: ProductDefinitionShape from StepRepr) returns FeaModel from StepFEA;
    FeaModel(me; PD: ProductDefinition from StepBasic) returns FeaModel from StepFEA;
    IdealShape(me; PD: ProductDefinition from StepBasic) returns ShapeRepresentation from StepShape;
    IdealShape(me; PDS: ProductDefinitionShape from StepRepr) returns ShapeRepresentation from StepShape;
   

--fields

end Construct;
