-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Loop from IGESSolid  inherits IGESEntity

        ---Purpose: defines Loop, Type <508> Form Number <1>
        --          in package IGESSolid
        --          A Loop entity specifies a bound of a face. It represents
        --          a connected collection of face boundaries, seams, and
        --          poles of a single face.
        --          
        --          From IGES-5.3, a Loop can be free with Form Number 0,
        --          else it is a bound of a face (it is the default)

uses

        HArray1OfIGESEntity                 from IGESData,
        HArray1OfInteger                    from TColStd,
        HArray1OfHArray1OfInteger           from IGESBasic,
        HArray1OfHArray1OfInteger_Handle    from IGESBasic,
        HArray1OfHArray1OfIGESEntity_Handle from IGESBasic

raises DimensionMismatch, OutOfRange

is

        Create returns mutable Loop;

        -- Specific Methods pertaining to the class

        Init (me                 : mutable;
              types              : HArray1OfInteger;
              edges              : HArray1OfIGESEntity;
              index              : HArray1OfInteger;
              orient             : HArray1OfInteger;
              nbParameterCurves  : HArray1OfInteger;
              isoparametricFlags : HArray1OfHArray1OfInteger_Handle;
              curves             : HArray1OfHArray1OfIGESEntity_Handle from
                                   IGESBasic)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class Loop
        --       - types              : 0 = Edge; 1 = Vertex
        --       - edges              : Pointer to the EdgeList or VertexList
        --       - index              : Index of the edge into the EdgeList
        --                              VertexList entity
        --       - orient             : Orientation flag of the edge
        --       - nbParameterCurves  : the number of parameter space curves
        --                              for each edge
        --       - isoparametricFlags : the isoparametric flag of the
        --                              parameter space curve
        --       - curves             : the parameter space curves
        -- raises exception if length of types, edges, index, orient and
        -- nbParameterCurves do not match or the length of
        -- isoparametricFlags and curves do not match

    	IsBound (me) returns Boolean;
	---Purpose : Tells if a Loop is a Bound (FN 1) else it is free (FN 0)

    	SetBound (me : mutable; bound : Boolean);
	---Purpose : Sets or Unset the Bound Status (from Form Number)
	--           Default is True

        NbEdges (me) returns Integer;
        ---Purpose : returns the number of edge tuples

        EdgeType (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : returns the type of Index'th edge (0 = Edge, 1 = Vertex)
        -- raises exception if Index <= 0 or Index > NbEdges()

        Edge (me; Index : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : return the EdgeList or VertexList corresponding to the Index
        -- raises exception if Index <= 0 or Index > NbEdges()

        Orientation (me; Index : Integer) returns Boolean
        raises OutOfRange;
        ---Purpose : returns the orientation flag corresponding to Index'th edge
        -- raises exception if Index <= 0 or Index > NbEdges()

        NbParameterCurves (me; Index : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : return the number of parameter space curves associated with
        -- Index'th Edge
        -- raises exception if Index <= 0 or Index > NbEdges()

        IsIsoparametric (me; EdgeIndex, CurveIndex : Integer)
            returns Boolean
        raises OutOfRange;
        -- returns the EdgeIndex'th edge's CurveIndex'th isoparametric flag
        -- raises exception if EdgeIndex <= 0 or EdgeIndex > NbEdges() or
        -- if CurveIndex <= 0 or CurveIndex > NbParameterCurves(EdgeIndex)

        ParametricCurve (me; EdgeIndex, CurveIndex : Integer) returns IGESEntity
        raises OutOfRange;
        ---Purpose : returns the CurveIndex'th parameter space curve associated with
        -- EdgeIndex'th edge
        -- raises exception if EdgeIndex <= 0 or EdgeIndex > NbEdges() or
        -- if CurveIndex <= 0 or CurveIndex > NbParameterCurves(EdgeIndex)

        ListIndex (me; num : Integer) returns Integer
        raises OutOfRange;
        ---Purpose : raises exception If num <= 0 or num > NbEdges()

fields

--
-- Class    : IGESSolid_Loop
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class Loop.
--
-- Reminder : A Loop instance is defined by :
--            either an edge, an orientation, and optional parameter
--            curves or (in case of a pole) a vertex and an optional
--            parameter space curve.
--

        theTypes              : HArray1OfInteger;
            -- array containing the type of the edge

        theEdges              : HArray1OfIGESEntity;
            -- array of Vertex List or Edge List entity

        theIndex              : HArray1OfInteger;
            -- array of list index into Vertex or Edge List entity

        theOrientationFlags   : HArray1OfInteger;
            -- array of orientation flags

        theNbParameterCurves  : HArray1OfInteger;
            -- no. of underlying parameter space curves

        theIsoparametricFlags : HArray1OfHArray1OfInteger_Handle;
            -- Isoparametric flags of the space curves

        theCurves             : HArray1OfHArray1OfIGESEntity_Handle
                                from IGESBasic;
            -- parameter space curves corresponding to the edges

end Loop;
