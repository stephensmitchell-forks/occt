-- File:	Unfolding_FunctionWithDerivative.cdl
-- Created:	Fri Sep  5 17:44:29 2008
-- Author:	Mikhail KLOKOV
--		<mkk@kurox>
---Copyright:	Open CASCADE 2008

class FunctionWithDerivative from Unfolding inherits FunctionWithDerivative from math
uses
    Array1OfXY from TColgp,
    Trsf2d from gp,
    Dir2d from gp
is

    Create (theMaster, theSlave: Array1OfXY from TColgp; 
    	    theDir: Dir2d from gp;
    	    theTrsf: Trsf2d from gp) 
    	returns FunctionWithDerivative from Unfolding;
    	---Purpose:

    Value(me: in out; X: Real; F: out Real)
        ---Purpose: Computes the value <F>of the function for the variable <X>.
    	--          Returns True if the calculation were successfully done, 
    	--          False otherwise.

    returns Boolean
    is redefined;
 
    Derivative(me: in out; X: Real; D: out Real)
        ---Purpose: Computes the derivative <D> of the function 
        --          for the variable <X>.
    	--           Returns True if the calculation were successfully done, 
    	--           False otherwise.

    returns Boolean
    is redefined;    

    Values(me: in out; X: Real; F, D: out Real)
    	---Purpose: Computes the value <F> and the derivative <D> of the 
    	--          function for the variable <X>.
    	--          Returns True if the calculation were successfully done,
    	--          False otherwise.

    returns Boolean
    is redefined;
    
    GetStateNumber (me: in out) returns Integer from Standard
    	is redefined;

    Area(me)
    	returns Real from Standard;
    
fields
    myMasterPolyLine: Array1OfXY from TColgp;
    mySlavePolyLine: Array1OfXY from TColgp;
    myTrsf: Trsf2d from gp;
    myShiftDir: Dir2d from gp;
    myShift: Real from Standard;
    myArea: Real from Standard;

end FunctionWithDerivative from Unfolding;
