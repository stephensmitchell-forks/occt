-- Created on: 1997-08-01
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package PCDM

uses

    CDM,TColStd,TCollection,Storage


is 
 
    enumeration ReaderStatus is  
	    RS_OK, 
	    RS_NoDriver, 
	    RS_UnknownFileDriver, 
	    RS_OpenError, 
	    RS_NoVersion, 
	    RS_NoSchema, 
	    RS_NoDocument, 
	    RS_ExtensionFailure,
	    RS_WrongStreamMode, 
	    RS_FormatFailure, 
	    RS_TypeFailure,
	    RS_TypeNotFoundInSchema, 
	    RS_UnrecognizedFileFormat, 
	    RS_MakeFailure,		     
	    RS_PermissionDenied, 
	    RS_DriverFailure,
	    RS_AlreadyRetrievedAndModified,
	    RS_AlreadyRetrieved,
	    RS_UnknownDocument,
	    RS_WrongResource,
	    RS_ReaderException,
	    RS_NoModel
    end ReaderStatus;
    
    enumeration StoreStatus is
	    SS_OK,
	    SS_DriverFailure,
	    SS_WriteFailure,
	    SS_Failure,
	    SS_Doc_IsNull,
	    SS_No_Obj,
	    SS_Info_Section_Error
    end StoreStatus;
    
    deferred class Document;
    class SequenceOfDocument instantiates Sequence from TCollection(Document from PCDM);

    deferred class Reader;
    deferred class Writer;
    deferred class RetrievalDriver;    
    deferred class StorageDriver;    

    class ReferenceIterator;    
---Category: exceptions

    exception DriverError inherits Failure from Standard;
    

    ---Category: classes for versioning  reading/writing og the headers.
    private class Reference;
    private class SequenceOfReference instantiates Sequence from TCollection(Reference from PCDM);
    private deferred class ReadWriter;
    private class ReadWriter_1;
    
    ---Category: type of FileDriver;
    --           
    private enumeration TypeOfFileDriver is TOFD_File, TOFD_CmpFile, TOFD_XmlFile, TOFD_Unknown
    end TypeOfFileDriver from PCDM;
    
    private pointer BaseDriverPointer to BaseDriver from Storage;    
    
---Category: drivers plugin.
--           
    FindStorageDriver(aDocument: Document from CDM) 
    returns Boolean from Standard;
    
    StorageDriver(aDocument: Document from CDM)
    returns StorageDriver from PCDM
    raises NoSuchObject from Standard;
    ---Purpose:   gets   in the  EuclidDesktop   resource  the plugin
    --          identifier of the driver plugs the driver.
    --          
    
    Schema(aSchemaName: ExtendedString from TCollection;
           anApplication: Application from CDM)
    ---Purpose: returns a schema to be used during a Store or Retrieve
    --          operation.
    --          Schema will plug the schema defined by
    --          the SchemaName method.
    returns Schema from Storage;
    
    FileDriverType(aFileName: AsciiString from TCollection; aBaseDriver: out BaseDriverPointer from PCDM)
    returns TypeOfFileDriver from PCDM
    is private;

    FileDriverType(theIStream: in out IStream from Standard; aBaseDriver: out BaseDriverPointer from PCDM)
    returns TypeOfFileDriver from PCDM
    is private;

end PCDM;
