-- Created on: 1991-02-21
-- Created by: Isabelle GRIGNON
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class   POnSurf from Extrema
    	---Purpose: Definition of a point on surface.

uses    Pnt from gp

is
    Create returns POnSurf;
    	---Purpose: Creation of an indefinite point on surface.
    	---C++: inline

    Create (U,V: Real; P: Pnt) returns POnSurf;
    	---Purpose: Creation of a point on surface with parameter 
    	--          values on the surface and a Pnt from gp.
    	---C++: inline

    Value (me) returns Pnt
    	---Purpose: Returns the 3d point.
    	---C++: return const&
    	---C++: inline
    	is static;

    Parameter (me; U,V: out Real) 
    	---Purpose: Returns the parameter values on the surface.
    	---C++: inline
    	is static;          
    
    Parameter (me : mutable; theU, theV: Real from Standard; theP : Pnt from gp) 
    	---Purpose: Sets the params of current POnSurf instance.
       --         (e.g. to the point to be projected).
    	---C++: inline
    	is static;          
    
    
fields
    myU: Real;
    myV: Real;
    myP: Pnt from gp;

end POnSurf;
